`timescale 1us/1ns
module Top ( A, B, C, D );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] D;
  wire   sign_A, sign_B, \two_en[1] , \expadd/N1 , \expadd/N2 , \expadd/N3 ,
         \expadd/N4 , \expadd/N5 , \expadd/N6 , \sub/N21 , \sub/N20 ,
         \sub/N19 , \sub/N18 , \sub/N17 , \sub/N16 , \sub/N15 , \sub/N14 ,
         \sub/N12 , \sub/N11 , \sub/N10 , \sub/N9 , \sub/N8 , \sub/N7 ,
         \sub/N6 , \sub/N5 , \selc/N209 , \selc/N208 , \selc/N207 ,
         \selc/N206 , \selc/N205 , \selc/N204 , \selc/N203 , \selc/N202 ,
         \selc/N201 , \selc/N200 , \selc/N199 , \selc/N198 , \selc/N197 ,
         \selc/N196 , \selc/N195 , \selc/N194 , \selc/N193 , \selc/N192 ,
         \selc/N191 , \selc/N190 , \selc/N189 , \selc/N188 , \selc/N187 ,
         \selc/N162 , \selc/N161 , \selc/N160 , \selc/N159 , \selc/N158 ,
         \selc/N157 , \selc/N156 , \selc/N155 , \selc/N154 , \selc/N153 ,
         \selc/N152 , \selc/N151 , \selc/N150 , \selc/N149 , \selc/N148 ,
         \selc/N147 , \selc/N146 , \selc/N145 , \selc/N144 , \selc/N143 ,
         \selc/N142 , \selc/N141 , \selc/N140 , \selc/N139 , \selc/N138 ,
         \selc/N137 , \selc/N136 , \selc/N135 , \selc/N134 , \selc/N133 ,
         \selc/N132 , \selc/N131 , \selc/N130 , \selc/N129 , \selc/N128 ,
         \selc/N127 , \selc/N126 , \selc/N125 , \selc/N124 , \selc/N123 ,
         \selc/N122 , \selc/N121 , \selc/N120 , \selc/N119 , \selc/N118 ,
         \selc/N117 , \selc/N116 , \selc/N115 , \selc/N114 , \align/N102 ,
         \align/N101 , \align/N100 , \align/N99 , \align/N98 , \align/N97 ,
         \align/N96 , \align/N95 , \align/N94 , \align/N93 , \align/N92 ,
         \align/N91 , \align/N90 , \align/N89 , \align/N88 , \align/N87 ,
         \align/N86 , \align/N85 , \align/N84 , \align/N83 , \align/N82 ,
         \align/N81 , \align/N80 , \align/N79 , \align/N78 , \align/N77 ,
         \align/N76 , \align/N75 , \align/N74 , \align/N73 , \align/N72 ,
         \align/N71 , \align/N70 , \align/N69 , \align/N68 , \align/N67 ,
         \align/N66 , \align/N65 , \align/N64 , \align/N63 , \align/N62 ,
         \align/N61 , \align/N60 , \align/N59 , \align/N58 , \align/N57 ,
         \align/N56 , \align/N55 , \align/N54 , \align/N52 , \align/N51 ,
         \align/N50 , \align/N49 , \align/N48 , \align/N47 , \align/N46 ,
         \align/N45 , \align/N44 , \align/N43 , \align/N42 , \align/N41 ,
         \align/N40 , \align/N39 , \align/N38 , \align/N37 , \align/N36 ,
         \align/N35 , \align/N34 , \align/N33 , \align/N32 , \align/N31 ,
         \align/N30 , \align/N29 , \align/N28 , \align/N27 , \align/N26 ,
         \align/N25 , \align/N24 , \align/N23 , \align/N22 , \align/N21 ,
         \align/N20 , \align/N19 , \align/N18 , \align/N17 , \align/N16 ,
         \align/N15 , \align/N14 , \align/N13 , \align/N12 , \align/N11 ,
         \align/N10 , \align/N9 , \align/N8 , \align/N7 , \align/N6 ,
         \align/N5 , \align/N4 , \sigadd/N51 , \sigadd/N50 , \sigadd/N49 ,
         \sigadd/N48 , \sigadd/N47 , \sigadd/N46 , \sigadd/N45 , \sigadd/N44 ,
         \sigadd/N43 , \sigadd/N42 , \sigadd/N41 , \sigadd/N40 , \sigadd/N39 ,
         \sigadd/N38 , \sigadd/N37 , \sigadd/N36 , \sigadd/N35 , \sigadd/N34 ,
         \sigadd/N33 , \sigadd/N32 , \sigadd/N31 , \sigadd/N30 , \sigadd/N29 ,
         \sigadd/N28 , \sigadd/N27 , \sigadd/N26 , \sigadd/N25 , \sigadd/N24 ,
         \sigadd/N23 , \sigadd/N22 , \sigadd/N21 , \sigadd/N20 , \sigadd/N19 ,
         \sigadd/N18 , \sigadd/N17 , \sigadd/N16 , \sigadd/N15 , \sigadd/N14 ,
         \sigadd/N13 , \sigadd/N12 , \sigadd/N11 , \sigadd/N10 , \sigadd/N9 ,
         \sigadd/N8 , \sigadd/N7 , \sigadd/N6 , \sigadd/N5 , \sigadd/N4 ,
         \sigadd/N3 , \sigadd/sig[0] , \sigadd/sig[1] , \sigadd/sig[2] ,
         \sigadd/sig[3] , \sigadd/sig[4] , \sigadd/n15 , \normal/N94 ,
         \normal/N91 , \normal/N90 , \normal/N89 , \normal/N88 , \normal/N79 ,
         \normal/N78 , \normal/N77 , \normal/N76 , \normal/N74 , \normal/N73 ,
         \normal/N72 , \normal/N71 , \normal/N70 , \normal/N69 , \normal/N68 ,
         \normal/N67 , \normal/N66 , \normal/N65 , \normal/N64 , \normal/N63 ,
         \normal/N62 , \normal/N61 , \normal/N60 , \normal/N59 , \normal/N58 ,
         \normal/N49 , \normal/N48 , \normal/N45 , \normal/N44 , \normal/N43 ,
         \normal/N42 , \normal/N33 , \normal/N32 , \normal/N31 , \normal/N30 ,
         \normal/N28 , \normal/N27 , \normal/N26 , \normal/N25 , \normal/N24 ,
         \normal/N23 , \normal/N22 , \normal/N15 , \normal/N14 , \normal/N11 ,
         \normal/N10 , \normal/N9 , \normal/N8 , \normal/N7 , \normal/N6 ,
         \normal/N5 , \normal/N4 , \normal/N3 , \normal/n30 , \normal/n29 ,
         \round/N30 , \round/N29 , \round/N28 , \round/N27 , \round/N26 ,
         \round/N25 , \round/N24 , \round/N23 , \round/N22 , \round/N21 ,
         \round/N20 , \round/N19 , \round/N18 , \round/N17 , \round/N16 ,
         \round/N15 , \round/N14 , \round/N13 , \round/N12 , \round/N11 ,
         \round/N10 , \round/N9 , \ctrl/N30 , \ctrl/N28 , \ctrl/N27 ,
         \ctrl/N14 , \ctrl/N12 , \ctrl/N11 , n39, \selc/r300/carry[45] ,
         \selc/r300/carry[44] , \selc/r300/carry[43] , \selc/r300/carry[42] ,
         \selc/r300/carry[41] , \selc/r300/carry[40] , \selc/r300/carry[39] ,
         \selc/r300/carry[38] , \selc/r300/carry[37] , \selc/r300/carry[36] ,
         \selc/r300/carry[35] , \selc/r300/carry[34] , \selc/r300/carry[33] ,
         \selc/r300/carry[32] , \selc/r300/carry[31] , \selc/r300/carry[30] ,
         \selc/r300/carry[29] , \selc/r300/carry[28] , \selc/r300/carry[27] ,
         \selc/r300/carry[26] , \selc/r300/carry[25] , \selc/r300/carry[24] ,
         \selc/r300/A[24] , \selc/r300/A[25] , \selc/r300/A[26] ,
         \selc/r300/A[27] , \selc/r300/A[28] , \selc/r300/A[29] ,
         \selc/r300/A[30] , \selc/r300/A[31] , \selc/r300/A[32] ,
         \selc/r300/A[33] , \selc/r300/A[34] , \selc/r300/A[35] ,
         \selc/r300/A[36] , \selc/r300/A[37] , \selc/r300/A[38] ,
         \selc/r300/A[39] , \selc/r300/A[40] , \selc/r300/A[41] ,
         \selc/r300/A[42] , \selc/r300/A[43] , \selc/r300/A[44] ,
         \selc/r300/A[45] , \align/sra_11/n757 , \align/sra_11/n754 ,
         \align/sra_11/n753 , \align/sra_11/n746 , \align/sra_11/n744 ,
         \align/sra_11/n743 , \align/sra_11/n742 , \align/sra_11/n741 ,
         \align/sra_11/n740 , \align/sra_11/n739 , \align/sra_11/n738 ,
         \align/sra_11/n737 , \align/sra_11/n736 , \align/sra_11/n735 ,
         \align/sra_11/n734 , \align/sra_11/n733 , \align/sra_11/n732 ,
         \align/sra_11/n731 , \align/sra_11/n730 , \align/sra_11/n729 ,
         \align/sra_11/n728 , \align/sra_11/n727 , \align/sra_11/n724 ,
         \align/sra_11/n723 , \align/sra_11/n722 , \align/sra_11/n721 ,
         \align/sra_11/n720 , \align/sra_11/n719 , \align/sra_11/n718 ,
         \align/sra_11/n717 , \align/sra_11/n716 , \align/sra_11/n715 ,
         \align/sra_11/n714 , \align/sra_11/n709 , \align/sra_11/n707 ,
         \align/sra_11/n706 , \align/sra_11/n705 , \align/sra_11/n704 ,
         \align/sra_11/n703 , \align/sra_11/n702 , \align/sra_11/n701 ,
         \align/sra_11/n700 , \align/sra_11/n699 , \align/sra_11/n698 ,
         \align/sra_11/n697 , \align/sra_11/n696 , \align/sra_11/n695 ,
         \align/sra_11/n694 , \align/sra_11/n693 , \align/sra_11/n690 ,
         \align/sra_11/n689 , \align/sra_11/n688 , \align/sra_11/n687 ,
         \align/sra_11/n686 , \align/sra_11/n685 , \align/sra_11/n684 ,
         \align/sra_11/n683 , \align/sra_11/n682 , \align/sra_11/n681 ,
         \align/sra_11/n678 , \align/sra_11/n677 , \align/sra_11/n676 ,
         \align/sra_11/n675 , \align/sra_11/n674 , \align/sra_11/n673 ,
         \align/sra_11/n672 , \align/sra_11/n671 , \align/sra_11/n670 ,
         \align/sra_11/n669 , \align/sra_11/n668 , \align/sra_11/n667 ,
         \align/sra_11/n666 , \align/sra_11/n665 , \align/sra_11/n664 ,
         \align/sra_11/n663 , \align/sra_11/n661 , \align/sra_11/n660 ,
         \align/sra_11/n659 , \align/sra_11/n658 , \align/sra_11/n657 ,
         \align/sra_11/n656 , \align/sra_11/n655 , \align/sra_11/n654 ,
         \align/sra_11/n653 , \align/sra_11/n652 , \align/sra_11/n651 ,
         \align/sra_11/n650 , \align/sra_11/n649 , \align/sra_11/n648 ,
         \align/sra_11/n647 , \align/sra_11/n646 , \align/sra_11/n645 ,
         \align/sra_11/n644 , \align/sra_11/n643 , \align/sra_11/n642 ,
         \align/sra_11/n636 , \align/sra_11/n634 , \align/sra_11/n633 ,
         \align/sra_11/n632 , \align/sra_11/n631 , \align/sra_11/n630 ,
         \align/sra_11/n629 , \align/sra_11/n628 , \align/sra_11/n627 ,
         \align/sra_11/n626 , \align/sra_11/n625 , \align/sra_11/n624 ,
         \align/sra_11/n623 , \align/sra_11/n622 , \align/sra_11/n621 ,
         \align/sra_11/n620 , \align/sra_11/n619 , \align/sra_11/n618 ,
         \align/sra_11/n617 , \align/sra_11/n616 , \align/sra_11/n615 ,
         \align/sra_11/n614 , \align/sra_11/n613 , \align/sra_11/n612 ,
         \align/sra_11/n611 , \align/sra_11/n610 , \align/sra_11/n609 ,
         \align/sra_11/n608 , \align/sra_11/n607 , \align/sra_11/n606 ,
         \align/sra_11/n605 , \align/sra_11/n604 , \align/sra_11/n603 ,
         \align/sra_11/n602 , \align/sra_11/n601 , \align/sra_11/n600 ,
         \align/sra_11/n599 , \align/sra_11/n598 , \align/sra_11/n597 ,
         \align/sra_11/n596 , \align/sra_11/n595 , \align/sra_11/n594 ,
         \align/sra_11/n593 , \align/sra_11/n592 , \align/sra_11/n591 ,
         \align/sra_11/n590 , \align/sra_11/n589 , \align/sra_11/n588 ,
         \align/sra_11/n587 , \align/sra_11/n586 , \align/sra_11/n585 ,
         \align/sra_11/n584 , \align/sra_11/n583 , \align/sra_11/n582 ,
         \align/sra_11/n581 , \align/sra_11/n573 , \align/sra_11/n571 ,
         \align/sra_11/n570 , \align/sra_11/n569 , \align/sra_11/n568 ,
         \align/sra_11/n567 , \align/sra_11/n566 , \align/sra_11/n565 ,
         \align/sra_11/n564 , \align/sra_11/n563 , \align/sra_11/n562 ,
         \align/sra_11/n561 , \align/sra_11/n560 , \align/sra_11/n559 ,
         \align/sra_11/n558 , \align/sra_11/n557 , \align/sra_11/n556 ,
         \align/sra_11/n555 , \align/sra_11/n554 , \align/sra_11/n553 ,
         \align/sra_11/n552 , \align/sra_11/n551 , \align/sra_11/n550 ,
         \align/sra_11/n549 , \align/sra_11/n548 , \align/sra_11/n547 ,
         \align/sra_11/n546 , \align/sra_11/n545 , \align/sra_11/n537 ,
         \align/sra_11/n535 , \align/sra_11/n534 , \align/sra_11/n533 ,
         \align/sra_11/n532 , \align/sra_11/n531 , \align/sra_11/n530 ,
         \align/sra_11/n529 , \align/sra_11/n528 , \align/sra_11/n527 ,
         \align/sra_11/n526 , \align/sra_11/n525 , \align/sra_11/n524 ,
         \align/sra_11/n523 , \align/sra_11/n522 , \align/sra_11/n521 ,
         \align/sra_11/n520 , \align/sra_11/n519 , \align/sra_11/n518 ,
         \align/sra_11/n517 , \align/sra_11/n516 , \align/sra_11/n515 ,
         \align/sra_11/n510 , \align/sra_11/n508 , \align/sra_11/n507 ,
         \align/sra_11/n506 , \align/sra_11/n501 , \align/sra_11/n499 ,
         \align/sra_11/n498 , \align/sra_11/n497 , \align/sra_11/n492 ,
         \align/sra_11/n490 , \align/sra_11/n489 , \align/sra_11/n488 ,
         \align/sra_11/n483 , \align/sra_11/n481 , \align/sra_11/n480 ,
         \align/sra_11/n479 , \align/sra_11/n478 , \align/sra_11/n476 ,
         \align/sra_11/n475 , \align/sra_11/n474 , \align/sra_11/n473 ,
         \align/sra_11/n472 , \align/sra_11/n471 , \align/sra_11/n469 ,
         \align/sra_11/n468 , \align/sra_11/n467 , \align/sra_11/n466 ,
         \align/sra_11/n465 , \align/sra_11/n464 , \align/sra_11/SH[1] ,
         \normal/srl_15/A[44] , \normal/srl_15/A[41] , \normal/srl_15/A[40] ,
         \normal/srl_15/A[36] , \normal/srl_15/A[32] , \normal/srl_15/A[29] ,
         \normal/srl_15/A[27] , \normal/srl_15/A[25] , \normal/srl_15/A[22] ,
         \normal/srl_15/A[21] , \normal/srl_15/A[12] , \normal/srl_15/A[11] ,
         \normal/srl_15/A[10] , \normal/srl_15/A[9] , \normal/srl_15/A[8] ,
         \normal/srl_15/A[6] , \normal/srl_15/A[4] , \normal/srl_15/A[1] ,
         \normal/srl_15/n248 , \normal/srl_15/n247 , \normal/srl_15/n246 ,
         \normal/srl_15/n245 , \normal/srl_15/n244 , \normal/srl_15/n243 ,
         \normal/srl_15/n242 , \normal/srl_15/n241 , \normal/srl_15/n240 ,
         \normal/srl_15/n239 , \normal/srl_15/n238 , \normal/srl_15/n237 ,
         \normal/srl_15/n236 , \normal/srl_15/n235 , \normal/srl_15/n234 ,
         \normal/srl_15/n233 , \normal/srl_15/n232 , \normal/srl_15/n231 ,
         \normal/srl_15/n230 , \normal/srl_15/n229 , \normal/srl_15/n228 ,
         \normal/srl_15/n227 , \normal/srl_15/n226 , \normal/srl_15/n225 ,
         \normal/srl_15/n224 , \normal/srl_15/n223 , \normal/srl_15/n222 ,
         \normal/srl_15/n221 , \normal/srl_15/n220 , \normal/srl_15/n219 ,
         \normal/srl_15/n218 , \normal/srl_15/n217 , \normal/srl_15/n216 ,
         \normal/srl_15/n215 , \normal/srl_15/n214 , \normal/srl_15/n213 ,
         \normal/srl_15/n212 , \normal/srl_15/n211 , \normal/srl_15/n210 ,
         \normal/srl_15/n209 , \normal/srl_15/n208 , \normal/srl_15/n207 ,
         \normal/srl_15/n206 , \normal/srl_15/n205 , \normal/srl_15/n204 ,
         \normal/srl_15/n203 , \normal/srl_15/n202 , \normal/srl_15/n201 ,
         \normal/srl_15/n200 , \normal/srl_15/n199 , \normal/srl_15/n198 ,
         \normal/srl_15/n197 , \normal/srl_15/n196 , \normal/srl_15/n195 ,
         \normal/srl_15/n194 , \normal/srl_15/n193 , \normal/srl_15/n192 ,
         \normal/srl_15/n191 , \normal/srl_15/n190 , \normal/srl_15/n189 ,
         \normal/srl_15/n188 , \normal/srl_15/n187 , \normal/srl_15/n186 ,
         \normal/srl_15/n185 , \normal/srl_15/n184 , \normal/srl_15/n183 ,
         \normal/srl_15/n182 , \normal/srl_15/n181 , \normal/srl_15/n175 ,
         \normal/srl_15/n174 , \normal/srl_15/n173 , \normal/srl_15/n169 ,
         \normal/srl_15/n166 , \normal/srl_15/n165 , \normal/srl_15/n164 ,
         \normal/srl_15/n163 , \normal/srl_15/n162 , \normal/srl_15/n161 ,
         \normal/srl_15/n160 , \normal/srl_15/n159 , \normal/srl_15/n158 ,
         \normal/srl_15/n157 , \normal/srl_15/n156 , \normal/srl_15/n155 ,
         \normal/srl_15/n154 , \normal/srl_15/n153 , \normal/srl_15/n152 ,
         \normal/srl_15/n151 , \normal/srl_15/n150 , \normal/srl_15/n149 ,
         \normal/srl_15/n148 , \normal/srl_15/n147 , \normal/srl_15/n146 ,
         \normal/srl_15/n145 , \normal/srl_15/n144 , \normal/srl_15/n143 ,
         \normal/srl_15/n142 , \normal/srl_15/n141 , \normal/srl_15/n140 ,
         \normal/srl_15/n139 , \normal/srl_15/n138 , \normal/srl_15/n137 ,
         \normal/srl_15/n136 , \normal/srl_15/n135 , \normal/srl_15/n134 ,
         \normal/srl_15/n133 , \normal/srl_15/n132 , \normal/srl_15/n131 ,
         \normal/srl_15/n130 , \normal/srl_15/n129 , \normal/srl_15/n128 ,
         \normal/srl_15/n127 , \normal/srl_15/n126 , \normal/srl_15/n125 ,
         \normal/srl_15/n124 , \normal/srl_15/n123 , \normal/srl_15/n122 ,
         \normal/srl_15/n121 , \normal/srl_15/n120 , \normal/srl_15/n119 ,
         \normal/srl_15/n118 , \normal/srl_15/n117 , \normal/srl_15/n116 ,
         \normal/srl_15/n115 , \normal/srl_15/n114 , \normal/srl_15/n113 ,
         \normal/srl_15/n112 , \normal/srl_15/n111 , \normal/srl_15/n110 ,
         \normal/srl_15/n109 , \normal/srl_15/n108 , \normal/srl_15/n107 ,
         \normal/srl_15/n106 , \normal/srl_15/n105 , \normal/srl_15/n104 ,
         \normal/srl_15/n103 , \normal/srl_15/n102 , \normal/srl_15/n101 ,
         \normal/srl_15/n100 , \normal/srl_15/n99 , \normal/srl_15/n98 ,
         \normal/srl_15/n97 , \normal/srl_15/n96 , \normal/srl_15/n95 ,
         \normal/srl_15/n94 , \normal/srl_15/n93 , \normal/srl_15/n92 ,
         \normal/srl_15/n91 , \normal/srl_15/n90 , \normal/srl_15/n89 ,
         \normal/srl_15/n88 , \normal/srl_15/n87 , \normal/srl_15/n86 ,
         \normal/srl_15/n85 , \normal/srl_15/n84 , \normal/srl_15/n83 ,
         \normal/srl_15/n82 , \normal/srl_15/n81 , \normal/srl_15/n80 ,
         \normal/srl_15/n79 , \normal/srl_15/n78 , \normal/srl_15/n77 ,
         \normal/srl_15/n76 , \normal/srl_15/n75 , \normal/srl_15/n74 ,
         \normal/srl_15/n73 , \normal/srl_15/n72 , \normal/srl_15/n71 ,
         \normal/srl_15/n70 , \normal/srl_15/n69 , \normal/srl_15/n68 ,
         \normal/srl_15/n67 , \normal/srl_15/n66 , \normal/srl_15/n65 ,
         \normal/srl_15/n64 , \normal/srl_15/n63 , \normal/srl_15/n62 ,
         \normal/srl_15/n61 , \normal/srl_15/n60 , \normal/srl_15/n59 ,
         \normal/srl_15/n58 , \normal/srl_15/n57 , \normal/srl_15/n56 ,
         \normal/srl_15/n55 , \normal/srl_15/n54 , \normal/srl_15/n53 ,
         \normal/srl_15/n52 , \normal/srl_15/n51 , \normal/srl_15/n50 ,
         \normal/srl_15/n49 , \normal/srl_15/n48 , \normal/srl_15/n47 ,
         \normal/srl_15/n46 , \normal/srl_15/n45 , \normal/srl_15/n44 ,
         \normal/srl_15/n43 , \normal/srl_15/n42 , \normal/srl_15/n41 ,
         \normal/srl_15/n40 , \normal/srl_15/n39 , \normal/srl_15/n38 ,
         \normal/srl_15/n37 , \normal/srl_15/n36 , \normal/srl_15/n35 ,
         \normal/srl_15/n34 , \normal/srl_15/n33 , \normal/srl_15/n32 ,
         \normal/srl_15/n31 , \normal/srl_15/n30 , \normal/srl_15/n29 ,
         \normal/srl_15/n28 , \normal/srl_15/n27 , \normal/srl_15/n26 ,
         \normal/srl_15/n25 , \normal/srl_15/n24 , \normal/srl_15/n23 ,
         \normal/srl_15/n22 , \normal/srl_15/n21 , \normal/srl_15/n20 ,
         \normal/srl_15/n19 , \normal/srl_15/n18 , \normal/srl_15/n17 ,
         \normal/srl_15/n16 , \normal/srl_15/n15 , \normal/srl_15/n14 ,
         \normal/srl_15/n13 , \normal/srl_15/n12 , \normal/srl_15/n11 ,
         \normal/srl_15/n10 , \normal/srl_15/n9 , \normal/srl_15/n8 ,
         \normal/srl_15/n7 , \normal/srl_15/n6 , \normal/srl_15/n5 ,
         \normal/srl_15/n4 , \normal/srl_15/n3 , \normal/srl_15/n2 ,
         \normal/srl_15/n1 , \ctrl/sub_0_root_add_0_root_sub_16/A[7] ,
         \ctrl/sub_0_root_add_0_root_sub_16/A[5] ,
         \ctrl/sub_0_root_add_0_root_sub_16/A[4] ,
         \ctrl/sub_0_root_add_0_root_sub_16/A[3] ,
         \ctrl/sub_0_root_add_0_root_sub_16/A[2] ,
         \ctrl/sub_0_root_add_0_root_sub_16/A[1] ,
         \ctrl/sub_0_root_add_0_root_sub_16/A[0] ,
         \ctrl/sub_0_root_add_0_root_sub_16/n40 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n38 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n36 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n35 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n34 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n33 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n32 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n31 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n29 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n27 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n26 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n25 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n24 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n23 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n21 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n19 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n14 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n12 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n10 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n8 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n7 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n6 ,
         \ctrl/sub_0_root_add_0_root_sub_16/n4 , \round/r298/n117 ,
         \round/r298/n116 , \round/r298/n113 , \round/r298/n112 ,
         \round/r298/n106 , \round/r298/n105 , \round/r298/n104 ,
         \round/r298/n103 , \round/r298/n95 , \round/r298/n87 ,
         \round/r298/n86 , \round/r298/n85 , \round/r298/n84 ,
         \round/r298/n83 , \round/r298/n81 , \round/r298/n80 ,
         \round/r298/n76 , \round/r298/n75 , \round/r298/n74 ,
         \round/r298/n73 , \round/r298/n70 , \round/r298/n69 ,
         \round/r298/n68 , \round/r298/n66 , \round/r298/n64 ,
         \round/r298/n63 , \round/r298/n62 , \round/r298/n61 ,
         \round/r298/n58 , \round/r298/n57 , \round/r298/n56 ,
         \round/r298/n53 , \round/r298/n52 , \round/r298/n51 ,
         \round/r298/n50 , \round/r298/n49 , \round/r298/n47 ,
         \round/r298/n46 , \round/r298/n45 , \round/r298/n44 ,
         \round/r298/n42 , \round/r298/n41 , \round/r298/n40 ,
         \round/r298/n36 , \round/r298/n35 , \round/r298/n31 ,
         \round/r298/n28 , \round/r298/n21 , \round/r298/n19 ,
         \round/r298/n18 , \round/r298/n17 , \round/r298/n16 , \round/r298/n9 ,
         \round/r298/n5 , \round/r298/n1 , \align/sra_10/n304 ,
         \align/sra_10/n303 , \align/sra_10/n302 , \align/sra_10/n301 ,
         \align/sra_10/n300 , \align/sra_10/n299 , \align/sra_10/n298 ,
         \align/sra_10/n297 , \align/sra_10/n296 , \align/sra_10/n295 ,
         \align/sra_10/n294 , \align/sra_10/n293 , \align/sra_10/n292 ,
         \align/sra_10/n291 , \align/sra_10/n290 , \align/sra_10/n289 ,
         \align/sra_10/n288 , \align/sra_10/n287 , \align/sra_10/n286 ,
         \align/sra_10/n285 , \align/sra_10/n284 , \align/sra_10/n283 ,
         \align/sra_10/n282 , \align/sra_10/n281 , \align/sra_10/n280 ,
         \align/sra_10/n279 , \align/sra_10/n278 , \align/sra_10/n277 ,
         \align/sra_10/n276 , \align/sra_10/n275 , \align/sra_10/n274 ,
         \align/sra_10/n273 , \align/sra_10/n272 , \align/sra_10/n271 ,
         \align/sra_10/n270 , \align/sra_10/n269 , \align/sra_10/n268 ,
         \align/sra_10/n267 , \align/sra_10/n266 , \align/sra_10/n265 ,
         \align/sra_10/n264 , \align/sra_10/n263 , \align/sra_10/n262 ,
         \align/sra_10/n261 , \align/sra_10/n260 , \align/sra_10/n259 ,
         \align/sra_10/n258 , \align/sra_10/n257 , \align/sra_10/n256 ,
         \align/sra_10/n255 , \align/sra_10/n254 , \align/sra_10/n250 ,
         \align/sra_10/n249 , \align/sra_10/n248 , \align/sra_10/n247 ,
         \align/sra_10/n246 , \align/sra_10/n245 , \align/sra_10/n244 ,
         \align/sra_10/n243 , \align/sra_10/n242 , \align/sra_10/n241 ,
         \align/sra_10/n240 , \align/sra_10/n239 , \align/sra_10/n238 ,
         \align/sra_10/n237 , \align/sra_10/n236 , \align/sra_10/n235 ,
         \align/sra_10/n234 , \align/sra_10/n233 , \align/sra_10/n232 ,
         \align/sra_10/n231 , \align/sra_10/n230 , \align/sra_10/n229 ,
         \align/sra_10/n228 , \align/sra_10/n227 , \align/sra_10/n226 ,
         \align/sra_10/n225 , \align/sra_10/n224 , \align/sra_10/n223 ,
         \align/sra_10/n222 , \align/sra_10/n221 , \align/sra_10/n220 ,
         \align/sra_10/n219 , \align/sra_10/n218 , \align/sra_10/n217 ,
         \align/sra_10/n216 , \align/sra_10/n215 , \align/sra_10/n214 ,
         \align/sra_10/n213 , \align/sra_10/n212 , \align/sra_10/n211 ,
         \align/sra_10/n210 , \align/sra_10/n209 , \align/sra_10/n208 ,
         \align/sra_10/n207 , \align/sra_10/n206 , \align/sra_10/n205 ,
         \align/sra_10/n204 , \align/sra_10/n203 , \align/sra_10/n202 ,
         \align/sra_10/n201 , \align/sra_10/n200 , \align/sra_10/n199 ,
         \align/sra_10/n198 , \align/sra_10/n197 , \align/sra_10/n196 ,
         \align/sra_10/n195 , \align/sra_10/n194 , \align/sra_10/n193 ,
         \align/sra_10/n192 , \align/sra_10/n191 , \align/sra_10/n190 ,
         \align/sra_10/n189 , \align/sra_10/n188 , \align/sra_10/n187 ,
         \align/sra_10/n186 , \align/sra_10/n185 , \align/sra_10/n184 ,
         \align/sra_10/n183 , \align/sra_10/n182 , \align/sra_10/n181 ,
         \align/sra_10/n180 , \align/sra_10/n179 , \align/sra_10/n178 ,
         \align/sra_10/n177 , \align/sra_10/n176 , \align/sra_10/n175 ,
         \align/sra_10/n174 , \align/sra_10/n173 , \align/sra_10/n172 ,
         \align/sra_10/n171 , \align/sra_10/n170 , \align/sra_10/n169 ,
         \align/sra_10/n168 , \align/sra_10/n167 , \align/sra_10/n166 ,
         \align/sra_10/n165 , \align/sra_10/n164 , \align/sra_10/n163 ,
         \align/sra_10/n162 , \align/sra_10/n161 , \align/sra_10/n160 ,
         \align/sra_10/n159 , \align/sra_10/n158 , \align/sra_10/n157 ,
         \align/sra_10/n156 , \align/sra_10/n155 , \align/sra_10/n154 ,
         \align/sra_10/n153 , \align/sra_10/n152 , \align/sra_10/n151 ,
         \align/sra_10/n150 , \align/sra_10/n149 , \align/sra_10/n148 ,
         \align/sra_10/n147 , \align/sra_10/n146 , \align/sra_10/n145 ,
         \align/sra_10/n144 , \align/sra_10/n143 , \align/sra_10/n142 ,
         \align/sra_10/n141 , \align/sra_10/n140 , \align/sra_10/n139 ,
         \align/sra_10/n138 , \align/sra_10/n137 , \align/sra_10/n136 ,
         \align/sra_10/n135 , \align/sra_10/n134 , \align/sra_10/n133 ,
         \align/sra_10/n132 , \align/sra_10/n131 , \align/sra_10/n130 ,
         \align/sra_10/n129 , \align/sra_10/n128 , \align/sra_10/n127 ,
         \align/sra_10/n126 , \align/sra_10/n125 , \align/sra_10/n124 ,
         \align/sra_10/n123 , \align/sra_10/n122 , \align/sra_10/n121 ,
         \align/sra_10/n120 , \align/sra_10/n119 , \align/sra_10/n118 ,
         \align/sra_10/n117 , \align/sra_10/n116 , \align/sra_10/n115 ,
         \align/sra_10/n114 , \align/sra_10/n113 , \align/sra_10/n112 ,
         \align/sra_10/n111 , \align/sra_10/n110 , \align/sra_10/n109 ,
         \align/sra_10/n108 , \align/sra_10/n107 , \align/sra_10/n106 ,
         \align/sra_10/n105 , \align/sra_10/n104 , \align/sra_10/n103 ,
         \align/sra_10/n102 , \align/sra_10/n101 , \align/sra_10/n100 ,
         \align/sra_10/n99 , \align/sra_10/n98 , \align/sra_10/n97 ,
         \align/sra_10/n96 , \align/sra_10/n95 , \align/sra_10/n94 ,
         \align/sra_10/n93 , \align/sra_10/n92 , \align/sra_10/n91 ,
         \align/sra_10/n90 , \align/sra_10/n89 , \align/sra_10/n88 ,
         \align/sra_10/n87 , \align/sra_10/n86 , \align/sra_10/n85 ,
         \align/sra_10/n84 , \align/sra_10/n83 , \align/sra_10/n82 ,
         \align/sra_10/n81 , \align/sra_10/n80 , \align/sra_10/n79 ,
         \align/sra_10/n78 , \align/sra_10/n77 , \align/sra_10/n76 ,
         \align/sra_10/n75 , \align/sra_10/n74 , \align/sra_10/n73 ,
         \align/sra_10/n72 , \align/sra_10/n71 , \align/sra_10/n70 ,
         \align/sra_10/n69 , \align/sra_10/n68 , \align/sra_10/n67 ,
         \align/sra_10/n66 , \align/sra_10/n65 , \align/sra_10/n64 ,
         \align/sra_10/n63 , \align/sra_10/n62 , \align/sra_10/n61 ,
         \align/sra_10/n60 , \align/sra_10/n59 , \align/sra_10/n58 ,
         \align/sra_10/n57 , \align/sra_10/n56 , \align/sra_10/n55 ,
         \align/sra_10/n54 , \align/sra_10/n53 , \align/sra_10/n52 ,
         \align/sra_10/n51 , \align/sra_10/n50 , \align/sra_10/n49 ,
         \align/sra_10/n48 , \align/sra_10/n47 , \align/sra_10/n46 ,
         \align/sra_10/n45 , \align/sra_10/n44 , \align/sra_10/n43 ,
         \align/sra_10/n42 , \align/sra_10/n41 , \align/sra_10/n40 ,
         \align/sra_10/n39 , \align/sra_10/n38 , \align/sra_10/n37 ,
         \align/sra_10/n36 , \align/sra_10/n35 , \align/sra_10/n34 ,
         \align/sra_10/n33 , \align/sra_10/n32 , \align/sra_10/n31 ,
         \align/sra_10/n30 , \align/sra_10/n29 , \align/sra_10/n28 ,
         \align/sra_10/n27 , \align/sra_10/n26 , \align/sra_10/n25 ,
         \align/sra_10/n24 , \align/sra_10/n23 , \align/sra_10/n22 ,
         \align/sra_10/n21 , \align/sra_10/n20 , \align/sra_10/n19 ,
         \align/sra_10/n18 , \align/sra_10/n17 , \align/sra_10/n16 ,
         \align/sra_10/n15 , \align/sra_10/n14 , \align/sra_10/n13 ,
         \align/sra_10/n12 , \align/sra_10/n11 , \align/sra_10/n10 ,
         \align/sra_10/n9 , \align/sra_10/n8 , \align/sra_10/n7 ,
         \align/sra_10/n6 , \align/sra_10/n5 , \align/sra_10/n4 ,
         \align/sra_10/n3 , \align/sra_10/n2 , \align/sra_10/n1 ,
         \normal/sll_15/n235 , \normal/sll_15/n234 , \normal/sll_15/n233 ,
         \normal/sll_15/n232 , \normal/sll_15/n231 , \normal/sll_15/n230 ,
         \normal/sll_15/n229 , \normal/sll_15/n228 , \normal/sll_15/n227 ,
         \normal/sll_15/n226 , \normal/sll_15/n225 , \normal/sll_15/n224 ,
         \normal/sll_15/n223 , \normal/sll_15/n222 , \normal/sll_15/n221 ,
         \normal/sll_15/n220 , \normal/sll_15/n219 , \normal/sll_15/n218 ,
         \normal/sll_15/n217 , \normal/sll_15/n216 , \normal/sll_15/n215 ,
         \normal/sll_15/n214 , \normal/sll_15/n213 , \normal/sll_15/n212 ,
         \normal/sll_15/n211 , \normal/sll_15/n210 , \normal/sll_15/n209 ,
         \normal/sll_15/n208 , \normal/sll_15/n207 , \normal/sll_15/n206 ,
         \normal/sll_15/n205 , \normal/sll_15/n204 , \normal/sll_15/n203 ,
         \normal/sll_15/n202 , \normal/sll_15/n201 , \normal/sll_15/n200 ,
         \normal/sll_15/n199 , \normal/sll_15/n198 , \normal/sll_15/n197 ,
         \normal/sll_15/n196 , \normal/sll_15/n195 , \normal/sll_15/n194 ,
         \normal/sll_15/n193 , \normal/sll_15/n192 , \normal/sll_15/n191 ,
         \normal/sll_15/n190 , \normal/sll_15/n189 , \normal/sll_15/n188 ,
         \normal/sll_15/n187 , \normal/sll_15/n186 , \normal/sll_15/n185 ,
         \normal/sll_15/n184 , \normal/sll_15/n183 , \normal/sll_15/n182 ,
         \normal/sll_15/n181 , \normal/sll_15/n180 , \normal/sll_15/n179 ,
         \normal/sll_15/n178 , \normal/sll_15/n177 , \normal/sll_15/n176 ,
         \normal/sll_15/n175 , \normal/sll_15/n174 , \normal/sll_15/n173 ,
         \normal/sll_15/n170 , \normal/sll_15/n169 , \normal/sll_15/n168 ,
         \normal/sll_15/n167 , \normal/sll_15/n158 , \normal/sll_15/n157 ,
         \normal/sll_15/n156 , \normal/sll_15/n155 , \normal/sll_15/n154 ,
         \normal/sll_15/n153 , \normal/sll_15/n152 , \normal/sll_15/n151 ,
         \normal/sll_15/n150 , \normal/sll_15/n149 , \normal/sll_15/n148 ,
         \normal/sll_15/n147 , \normal/sll_15/n146 , \normal/sll_15/n145 ,
         \normal/sll_15/n144 , \normal/sll_15/n143 , \normal/sll_15/n142 ,
         \normal/sll_15/n141 , \normal/sll_15/n140 , \normal/sll_15/n139 ,
         \normal/sll_15/n138 , \normal/sll_15/n137 , \normal/sll_15/n136 ,
         \normal/sll_15/n135 , \normal/sll_15/n134 , \normal/sll_15/n133 ,
         \normal/sll_15/n132 , \normal/sll_15/n131 , \normal/sll_15/n130 ,
         \normal/sll_15/n129 , \normal/sll_15/n128 , \normal/sll_15/n127 ,
         \normal/sll_15/n126 , \normal/sll_15/n125 , \normal/sll_15/n124 ,
         \normal/sll_15/n123 , \normal/sll_15/n122 , \normal/sll_15/n121 ,
         \normal/sll_15/n120 , \normal/sll_15/n119 , \normal/sll_15/n118 ,
         \normal/sll_15/n117 , \normal/sll_15/n116 , \normal/sll_15/n115 ,
         \normal/sll_15/n114 , \normal/sll_15/n113 , \normal/sll_15/n112 ,
         \normal/sll_15/n111 , \normal/sll_15/n110 , \normal/sll_15/n109 ,
         \normal/sll_15/n108 , \normal/sll_15/n107 , \normal/sll_15/n106 ,
         \normal/sll_15/n105 , \normal/sll_15/n104 , \normal/sll_15/n103 ,
         \normal/sll_15/n102 , \normal/sll_15/n101 , \normal/sll_15/n100 ,
         \normal/sll_15/n99 , \normal/sll_15/n98 , \normal/sll_15/n97 ,
         \normal/sll_15/n96 , \normal/sll_15/n95 , \normal/sll_15/n94 ,
         \normal/sll_15/n93 , \normal/sll_15/n92 , \normal/sll_15/n91 ,
         \normal/sll_15/n90 , \normal/sll_15/n89 , \normal/sll_15/n88 ,
         \normal/sll_15/n87 , \normal/sll_15/n86 , \normal/sll_15/n85 ,
         \normal/sll_15/n84 , \normal/sll_15/n83 , \normal/sll_15/n82 ,
         \normal/sll_15/n81 , \normal/sll_15/n80 , \normal/sll_15/n79 ,
         \normal/sll_15/n78 , \normal/sll_15/n77 , \normal/sll_15/n76 ,
         \normal/sll_15/n75 , \normal/sll_15/n74 , \normal/sll_15/n73 ,
         \normal/sll_15/n72 , \normal/sll_15/n71 , \normal/sll_15/n70 ,
         \normal/sll_15/n69 , \normal/sll_15/n68 , \normal/sll_15/n67 ,
         \normal/sll_15/n66 , \normal/sll_15/n65 , \normal/sll_15/n64 ,
         \normal/sll_15/n63 , \normal/sll_15/n62 , \normal/sll_15/n61 ,
         \normal/sll_15/n60 , \normal/sll_15/n59 , \normal/sll_15/n58 ,
         \normal/sll_15/n57 , \normal/sll_15/n56 , \normal/sll_15/n55 ,
         \normal/sll_15/n54 , \normal/sll_15/n53 , \normal/sll_15/n52 ,
         \normal/sll_15/n51 , \normal/sll_15/n50 , \normal/sll_15/n49 ,
         \normal/sll_15/n48 , \normal/sll_15/n47 , \normal/sll_15/n46 ,
         \normal/sll_15/n45 , \normal/sll_15/n44 , \normal/sll_15/n43 ,
         \normal/sll_15/n42 , \normal/sll_15/n41 , \normal/sll_15/n40 ,
         \normal/sll_15/n39 , \normal/sll_15/n38 , \normal/sll_15/n37 ,
         \normal/sll_15/n36 , \normal/sll_15/n35 , \normal/sll_15/n34 ,
         \normal/sll_15/n33 , \normal/sll_15/n32 , \normal/sll_15/n31 ,
         \normal/sll_15/n30 , \normal/sll_15/n29 , \normal/sll_15/n28 ,
         \normal/sll_15/n27 , \normal/sll_15/n26 , \normal/sll_15/n25 ,
         \normal/sll_15/n24 , \normal/sll_15/n23 , \normal/sll_15/n22 ,
         \normal/sll_15/n21 , \normal/sll_15/n20 , \normal/sll_15/n19 ,
         \normal/sll_15/n18 , \normal/sll_15/n17 , \normal/sll_15/n16 ,
         \normal/sll_15/n15 , \normal/sll_15/n14 , \normal/sll_15/n13 ,
         \normal/sll_15/n12 , \normal/sll_15/n11 , \normal/sll_15/n10 ,
         \normal/sll_15/n9 , \normal/sll_15/n5 , \normal/sll_15/n1 ,
         \ctrl/add_1_root_add_16_2/A[4] , \ctrl/add_1_root_add_16_2/A[2] ,
         \ctrl/add_1_root_add_16_2/A[0] , \ctrl/add_1_root_add_16_2/n67 ,
         \ctrl/add_1_root_add_16_2/n65 , \ctrl/add_1_root_add_16_2/n62 ,
         \ctrl/add_1_root_add_16_2/n60 , \ctrl/add_1_root_add_16_2/n58 ,
         \ctrl/add_1_root_add_16_2/n57 , \ctrl/add_1_root_add_16_2/n49 ,
         \ctrl/add_1_root_add_16_2/n48 , \ctrl/add_1_root_add_16_2/n44 ,
         \ctrl/add_1_root_add_16_2/n41 , \ctrl/add_1_root_add_16_2/n40 ,
         \ctrl/add_1_root_add_16_2/n39 , \ctrl/add_1_root_add_16_2/n38 ,
         \ctrl/add_1_root_add_16_2/n37 , \ctrl/add_1_root_add_16_2/n36 ,
         \ctrl/add_1_root_add_16_2/n31 , \ctrl/add_1_root_add_16_2/n30 ,
         \ctrl/add_1_root_add_16_2/n28 , \ctrl/add_1_root_add_16_2/n26 ,
         \ctrl/add_1_root_add_16_2/n24 , \ctrl/add_1_root_add_16_2/n23 ,
         \ctrl/add_1_root_add_16_2/n22 , \ctrl/add_1_root_add_16_2/n21 ,
         \ctrl/add_1_root_add_16_2/n19 , \ctrl/add_1_root_add_16_2/n18 ,
         \ctrl/add_1_root_add_16_2/n17 , \ctrl/add_1_root_add_16_2/n16 ,
         \ctrl/add_1_root_add_16_2/n15 , \ctrl/add_1_root_add_16_2/n13 ,
         \ctrl/add_1_root_add_16_2/n8 , \ctrl/add_1_root_add_16_2/n7 ,
         \ctrl/add_1_root_add_16_2/n6 , \ctrl/add_1_root_add_16_2/n5 ,
         \ctrl/add_1_root_add_16_2/n3 , \mul/mult_6/n1459 , \mul/mult_6/n1458 ,
         \mul/mult_6/n1457 , \mul/mult_6/n1456 , \mul/mult_6/n1455 ,
         \mul/mult_6/n1454 , \mul/mult_6/n1453 , \mul/mult_6/n1452 ,
         \mul/mult_6/n1451 , \mul/mult_6/n1450 , \mul/mult_6/n1449 ,
         \mul/mult_6/n1448 , \mul/mult_6/n1447 , \mul/mult_6/n1446 ,
         \mul/mult_6/n1445 , \mul/mult_6/n1444 , \mul/mult_6/n1443 ,
         \mul/mult_6/n1442 , \mul/mult_6/n1441 , \mul/mult_6/n1440 ,
         \mul/mult_6/n1439 , \mul/mult_6/n1438 , \mul/mult_6/n1437 ,
         \mul/mult_6/n1436 , \mul/mult_6/n1411 , \mul/mult_6/n1408 ,
         \mul/mult_6/n1407 , \mul/mult_6/n1405 , \mul/mult_6/n1402 ,
         \mul/mult_6/n1400 , \mul/mult_6/n1398 , \mul/mult_6/n1396 ,
         \mul/mult_6/n1394 , \mul/mult_6/n1392 , \mul/mult_6/n1391 ,
         \mul/mult_6/n1390 , \mul/mult_6/n1387 , \mul/mult_6/n1386 ,
         \mul/mult_6/n1383 , \mul/mult_6/n1382 , \mul/mult_6/n1380 ,
         \mul/mult_6/n1377 , \mul/mult_6/n1375 , \mul/mult_6/n1373 ,
         \mul/mult_6/n1371 , \mul/mult_6/n1369 , \mul/mult_6/n1367 ,
         \mul/mult_6/n1366 , \mul/mult_6/n1365 , \mul/mult_6/n1364 ,
         \mul/mult_6/n1363 , \mul/mult_6/n1360 , \mul/mult_6/n1359 ,
         \mul/mult_6/n1358 , \mul/mult_6/n1357 , \mul/mult_6/n1356 ,
         \mul/mult_6/n1355 , \mul/mult_6/n1354 , \mul/mult_6/n1353 ,
         \mul/mult_6/n1352 , \mul/mult_6/n1351 , \mul/mult_6/n1350 ,
         \mul/mult_6/n1349 , \mul/mult_6/n1348 , \mul/mult_6/n1347 ,
         \mul/mult_6/n1346 , \mul/mult_6/n1345 , \mul/mult_6/n1344 ,
         \mul/mult_6/n1343 , \mul/mult_6/n1342 , \mul/mult_6/n1341 ,
         \mul/mult_6/n1340 , \mul/mult_6/n1339 , \mul/mult_6/n1338 ,
         \mul/mult_6/n1336 , \mul/mult_6/n1335 , \mul/mult_6/n1334 ,
         \mul/mult_6/n1333 , \mul/mult_6/n1332 , \mul/mult_6/n1331 ,
         \mul/mult_6/n1330 , \mul/mult_6/n1329 , \mul/mult_6/n1328 ,
         \mul/mult_6/n1327 , \mul/mult_6/n1326 , \mul/mult_6/n1325 ,
         \mul/mult_6/n1324 , \mul/mult_6/n1323 , \mul/mult_6/n1322 ,
         \mul/mult_6/n1321 , \mul/mult_6/n1320 , \mul/mult_6/n1319 ,
         \mul/mult_6/n1318 , \mul/mult_6/n1317 , \mul/mult_6/n1316 ,
         \mul/mult_6/n1315 , \mul/mult_6/n1314 , \mul/mult_6/n1313 ,
         \mul/mult_6/n1312 , \mul/mult_6/n1311 , \mul/mult_6/n1308 ,
         \mul/mult_6/n1307 , \mul/mult_6/n1306 , \mul/mult_6/n1305 ,
         \mul/mult_6/n1304 , \mul/mult_6/n1303 , \mul/mult_6/n1302 ,
         \mul/mult_6/n1301 , \mul/mult_6/n1300 , \mul/mult_6/n1299 ,
         \mul/mult_6/n1298 , \mul/mult_6/n1297 , \mul/mult_6/n1296 ,
         \mul/mult_6/n1295 , \mul/mult_6/n1294 , \mul/mult_6/n1293 ,
         \mul/mult_6/n1292 , \mul/mult_6/n1291 , \mul/mult_6/n1290 ,
         \mul/mult_6/n1289 , \mul/mult_6/n1288 , \mul/mult_6/n1287 ,
         \mul/mult_6/n1286 , \mul/mult_6/n1284 , \mul/mult_6/n1283 ,
         \mul/mult_6/n1282 , \mul/mult_6/n1281 , \mul/mult_6/n1280 ,
         \mul/mult_6/n1279 , \mul/mult_6/n1278 , \mul/mult_6/n1277 ,
         \mul/mult_6/n1276 , \mul/mult_6/n1275 , \mul/mult_6/n1274 ,
         \mul/mult_6/n1273 , \mul/mult_6/n1272 , \mul/mult_6/n1271 ,
         \mul/mult_6/n1270 , \mul/mult_6/n1269 , \mul/mult_6/n1268 ,
         \mul/mult_6/n1267 , \mul/mult_6/n1266 , \mul/mult_6/n1265 ,
         \mul/mult_6/n1264 , \mul/mult_6/n1263 , \mul/mult_6/n1262 ,
         \mul/mult_6/n1261 , \mul/mult_6/n1260 , \mul/mult_6/n1259 ,
         \mul/mult_6/n1256 , \mul/mult_6/n1255 , \mul/mult_6/n1254 ,
         \mul/mult_6/n1253 , \mul/mult_6/n1252 , \mul/mult_6/n1251 ,
         \mul/mult_6/n1250 , \mul/mult_6/n1249 , \mul/mult_6/n1248 ,
         \mul/mult_6/n1247 , \mul/mult_6/n1246 , \mul/mult_6/n1245 ,
         \mul/mult_6/n1244 , \mul/mult_6/n1243 , \mul/mult_6/n1242 ,
         \mul/mult_6/n1241 , \mul/mult_6/n1240 , \mul/mult_6/n1239 ,
         \mul/mult_6/n1238 , \mul/mult_6/n1237 , \mul/mult_6/n1236 ,
         \mul/mult_6/n1235 , \mul/mult_6/n1234 , \mul/mult_6/n1232 ,
         \mul/mult_6/n1231 , \mul/mult_6/n1230 , \mul/mult_6/n1229 ,
         \mul/mult_6/n1228 , \mul/mult_6/n1227 , \mul/mult_6/n1226 ,
         \mul/mult_6/n1225 , \mul/mult_6/n1224 , \mul/mult_6/n1223 ,
         \mul/mult_6/n1222 , \mul/mult_6/n1221 , \mul/mult_6/n1220 ,
         \mul/mult_6/n1219 , \mul/mult_6/n1218 , \mul/mult_6/n1217 ,
         \mul/mult_6/n1216 , \mul/mult_6/n1215 , \mul/mult_6/n1214 ,
         \mul/mult_6/n1213 , \mul/mult_6/n1212 , \mul/mult_6/n1211 ,
         \mul/mult_6/n1210 , \mul/mult_6/n1209 , \mul/mult_6/n1208 ,
         \mul/mult_6/n1207 , \mul/mult_6/n1204 , \mul/mult_6/n1203 ,
         \mul/mult_6/n1202 , \mul/mult_6/n1201 , \mul/mult_6/n1200 ,
         \mul/mult_6/n1199 , \mul/mult_6/n1198 , \mul/mult_6/n1197 ,
         \mul/mult_6/n1196 , \mul/mult_6/n1195 , \mul/mult_6/n1194 ,
         \mul/mult_6/n1193 , \mul/mult_6/n1192 , \mul/mult_6/n1191 ,
         \mul/mult_6/n1190 , \mul/mult_6/n1189 , \mul/mult_6/n1188 ,
         \mul/mult_6/n1187 , \mul/mult_6/n1186 , \mul/mult_6/n1185 ,
         \mul/mult_6/n1184 , \mul/mult_6/n1183 , \mul/mult_6/n1182 ,
         \mul/mult_6/n1180 , \mul/mult_6/n1179 , \mul/mult_6/n1178 ,
         \mul/mult_6/n1177 , \mul/mult_6/n1176 , \mul/mult_6/n1175 ,
         \mul/mult_6/n1174 , \mul/mult_6/n1173 , \mul/mult_6/n1172 ,
         \mul/mult_6/n1171 , \mul/mult_6/n1170 , \mul/mult_6/n1169 ,
         \mul/mult_6/n1168 , \mul/mult_6/n1167 , \mul/mult_6/n1166 ,
         \mul/mult_6/n1165 , \mul/mult_6/n1164 , \mul/mult_6/n1163 ,
         \mul/mult_6/n1162 , \mul/mult_6/n1161 , \mul/mult_6/n1160 ,
         \mul/mult_6/n1159 , \mul/mult_6/n1158 , \mul/mult_6/n1157 ,
         \mul/mult_6/n1156 , \mul/mult_6/n1155 , \mul/mult_6/n1152 ,
         \mul/mult_6/n1151 , \mul/mult_6/n1150 , \mul/mult_6/n1149 ,
         \mul/mult_6/n1148 , \mul/mult_6/n1147 , \mul/mult_6/n1146 ,
         \mul/mult_6/n1145 , \mul/mult_6/n1144 , \mul/mult_6/n1143 ,
         \mul/mult_6/n1142 , \mul/mult_6/n1141 , \mul/mult_6/n1140 ,
         \mul/mult_6/n1139 , \mul/mult_6/n1138 , \mul/mult_6/n1137 ,
         \mul/mult_6/n1136 , \mul/mult_6/n1135 , \mul/mult_6/n1134 ,
         \mul/mult_6/n1133 , \mul/mult_6/n1132 , \mul/mult_6/n1131 ,
         \mul/mult_6/n1130 , \mul/mult_6/n1128 , \mul/mult_6/n1127 ,
         \mul/mult_6/n1126 , \mul/mult_6/n1125 , \mul/mult_6/n1124 ,
         \mul/mult_6/n1123 , \mul/mult_6/n1122 , \mul/mult_6/n1121 ,
         \mul/mult_6/n1120 , \mul/mult_6/n1119 , \mul/mult_6/n1118 ,
         \mul/mult_6/n1117 , \mul/mult_6/n1116 , \mul/mult_6/n1115 ,
         \mul/mult_6/n1114 , \mul/mult_6/n1113 , \mul/mult_6/n1112 ,
         \mul/mult_6/n1111 , \mul/mult_6/n1110 , \mul/mult_6/n1109 ,
         \mul/mult_6/n1108 , \mul/mult_6/n1107 , \mul/mult_6/n1106 ,
         \mul/mult_6/n1105 , \mul/mult_6/n1104 , \mul/mult_6/n1103 ,
         \mul/mult_6/n1100 , \mul/mult_6/n1099 , \mul/mult_6/n1098 ,
         \mul/mult_6/n1097 , \mul/mult_6/n1096 , \mul/mult_6/n1095 ,
         \mul/mult_6/n1094 , \mul/mult_6/n1093 , \mul/mult_6/n1092 ,
         \mul/mult_6/n1091 , \mul/mult_6/n1090 , \mul/mult_6/n1089 ,
         \mul/mult_6/n1088 , \mul/mult_6/n1087 , \mul/mult_6/n1086 ,
         \mul/mult_6/n1085 , \mul/mult_6/n1084 , \mul/mult_6/n1083 ,
         \mul/mult_6/n1082 , \mul/mult_6/n1081 , \mul/mult_6/n1080 ,
         \mul/mult_6/n1079 , \mul/mult_6/n1078 , \mul/mult_6/n1076 ,
         \mul/mult_6/n1075 , \mul/mult_6/n1074 , \mul/mult_6/n1073 ,
         \mul/mult_6/n1072 , \mul/mult_6/n1071 , \mul/mult_6/n1070 ,
         \mul/mult_6/n1069 , \mul/mult_6/n1068 , \mul/mult_6/n1067 ,
         \mul/mult_6/n1066 , \mul/mult_6/n1065 , \mul/mult_6/n1064 ,
         \mul/mult_6/n1063 , \mul/mult_6/n1062 , \mul/mult_6/n1061 ,
         \mul/mult_6/n1060 , \mul/mult_6/n1059 , \mul/mult_6/n1058 ,
         \mul/mult_6/n1057 , \mul/mult_6/n1056 , \mul/mult_6/n1055 ,
         \mul/mult_6/n1054 , \mul/mult_6/n1053 , \mul/mult_6/n1052 ,
         \mul/mult_6/n1051 , \mul/mult_6/n1048 , \mul/mult_6/n1047 ,
         \mul/mult_6/n1046 , \mul/mult_6/n1045 , \mul/mult_6/n1044 ,
         \mul/mult_6/n1043 , \mul/mult_6/n1042 , \mul/mult_6/n1041 ,
         \mul/mult_6/n1040 , \mul/mult_6/n1039 , \mul/mult_6/n1038 ,
         \mul/mult_6/n1037 , \mul/mult_6/n1036 , \mul/mult_6/n1035 ,
         \mul/mult_6/n1034 , \mul/mult_6/n1033 , \mul/mult_6/n1032 ,
         \mul/mult_6/n1031 , \mul/mult_6/n1030 , \mul/mult_6/n1029 ,
         \mul/mult_6/n1028 , \mul/mult_6/n1027 , \mul/mult_6/n1026 ,
         \mul/mult_6/n1024 , \mul/mult_6/n1023 , \mul/mult_6/n1022 ,
         \mul/mult_6/n1021 , \mul/mult_6/n1020 , \mul/mult_6/n1019 ,
         \mul/mult_6/n1018 , \mul/mult_6/n1017 , \mul/mult_6/n1016 ,
         \mul/mult_6/n1015 , \mul/mult_6/n1014 , \mul/mult_6/n1013 ,
         \mul/mult_6/n1012 , \mul/mult_6/n1011 , \mul/mult_6/n1010 ,
         \mul/mult_6/n1009 , \mul/mult_6/n1008 , \mul/mult_6/n1007 ,
         \mul/mult_6/n1006 , \mul/mult_6/n1005 , \mul/mult_6/n1004 ,
         \mul/mult_6/n1003 , \mul/mult_6/n1002 , \mul/mult_6/n1001 ,
         \mul/mult_6/n1000 , \mul/mult_6/n999 , \mul/mult_6/n996 ,
         \mul/mult_6/n995 , \mul/mult_6/n994 , \mul/mult_6/n993 ,
         \mul/mult_6/n992 , \mul/mult_6/n991 , \mul/mult_6/n990 ,
         \mul/mult_6/n989 , \mul/mult_6/n988 , \mul/mult_6/n987 ,
         \mul/mult_6/n986 , \mul/mult_6/n985 , \mul/mult_6/n984 ,
         \mul/mult_6/n983 , \mul/mult_6/n982 , \mul/mult_6/n981 ,
         \mul/mult_6/n980 , \mul/mult_6/n979 , \mul/mult_6/n978 ,
         \mul/mult_6/n977 , \mul/mult_6/n976 , \mul/mult_6/n975 ,
         \mul/mult_6/n974 , \mul/mult_6/n946 , \mul/mult_6/n945 ,
         \mul/mult_6/n944 , \mul/mult_6/n943 , \mul/mult_6/n942 ,
         \mul/mult_6/n941 , \mul/mult_6/n940 , \mul/mult_6/n939 ,
         \mul/mult_6/n938 , \mul/mult_6/n937 , \mul/mult_6/n936 ,
         \mul/mult_6/n935 , \mul/mult_6/n934 , \mul/mult_6/n933 ,
         \mul/mult_6/n932 , \mul/mult_6/n931 , \mul/mult_6/n930 ,
         \mul/mult_6/n929 , \mul/mult_6/n928 , \mul/mult_6/n927 ,
         \mul/mult_6/n926 , \mul/mult_6/n925 , \mul/mult_6/n924 ,
         \mul/mult_6/n923 , \mul/mult_6/n922 , \mul/mult_6/n921 ,
         \mul/mult_6/n919 , \mul/mult_6/n918 , \mul/mult_6/n917 ,
         \mul/mult_6/n916 , \mul/mult_6/n915 , \mul/mult_6/n914 ,
         \mul/mult_6/n913 , \mul/mult_6/n912 , \mul/mult_6/n911 ,
         \mul/mult_6/n910 , \mul/mult_6/n909 , \mul/mult_6/n908 ,
         \mul/mult_6/n907 , \mul/mult_6/n906 , \mul/mult_6/n905 ,
         \mul/mult_6/n904 , \mul/mult_6/n903 , \mul/mult_6/n902 ,
         \mul/mult_6/n901 , \mul/mult_6/n900 , \mul/mult_6/n899 ,
         \mul/mult_6/n898 , \mul/mult_6/n897 , \mul/mult_6/n896 ,
         \mul/mult_6/n895 , \mul/mult_6/n894 , \mul/mult_6/n892 ,
         \mul/mult_6/n891 , \mul/mult_6/n890 , \mul/mult_6/n889 ,
         \mul/mult_6/n888 , \mul/mult_6/n887 , \mul/mult_6/n886 ,
         \mul/mult_6/n885 , \mul/mult_6/n884 , \mul/mult_6/n883 ,
         \mul/mult_6/n882 , \mul/mult_6/n881 , \mul/mult_6/n880 ,
         \mul/mult_6/n879 , \mul/mult_6/n878 , \mul/mult_6/n877 ,
         \mul/mult_6/n876 , \mul/mult_6/n875 , \mul/mult_6/n874 ,
         \mul/mult_6/n873 , \mul/mult_6/n872 , \mul/mult_6/n871 ,
         \mul/mult_6/n870 , \mul/mult_6/n869 , \mul/mult_6/n868 ,
         \mul/mult_6/n867 , \mul/mult_6/n865 , \mul/mult_6/n864 ,
         \mul/mult_6/n863 , \mul/mult_6/n862 , \mul/mult_6/n861 ,
         \mul/mult_6/n860 , \mul/mult_6/n859 , \mul/mult_6/n858 ,
         \mul/mult_6/n857 , \mul/mult_6/n856 , \mul/mult_6/n855 ,
         \mul/mult_6/n854 , \mul/mult_6/n853 , \mul/mult_6/n852 ,
         \mul/mult_6/n851 , \mul/mult_6/n850 , \mul/mult_6/n849 ,
         \mul/mult_6/n848 , \mul/mult_6/n847 , \mul/mult_6/n846 ,
         \mul/mult_6/n845 , \mul/mult_6/n844 , \mul/mult_6/n843 ,
         \mul/mult_6/n842 , \mul/mult_6/n841 , \mul/mult_6/n840 ,
         \mul/mult_6/n838 , \mul/mult_6/n837 , \mul/mult_6/n836 ,
         \mul/mult_6/n835 , \mul/mult_6/n834 , \mul/mult_6/n833 ,
         \mul/mult_6/n832 , \mul/mult_6/n831 , \mul/mult_6/n830 ,
         \mul/mult_6/n829 , \mul/mult_6/n828 , \mul/mult_6/n827 ,
         \mul/mult_6/n826 , \mul/mult_6/n825 , \mul/mult_6/n824 ,
         \mul/mult_6/n823 , \mul/mult_6/n822 , \mul/mult_6/n821 ,
         \mul/mult_6/n820 , \mul/mult_6/n819 , \mul/mult_6/n818 ,
         \mul/mult_6/n817 , \mul/mult_6/n816 , \mul/mult_6/n815 ,
         \mul/mult_6/n814 , \mul/mult_6/n813 , \mul/mult_6/n811 ,
         \mul/mult_6/n810 , \mul/mult_6/n809 , \mul/mult_6/n808 ,
         \mul/mult_6/n807 , \mul/mult_6/n806 , \mul/mult_6/n805 ,
         \mul/mult_6/n804 , \mul/mult_6/n803 , \mul/mult_6/n802 ,
         \mul/mult_6/n801 , \mul/mult_6/n800 , \mul/mult_6/n799 ,
         \mul/mult_6/n798 , \mul/mult_6/n797 , \mul/mult_6/n796 ,
         \mul/mult_6/n795 , \mul/mult_6/n794 , \mul/mult_6/n793 ,
         \mul/mult_6/n792 , \mul/mult_6/n791 , \mul/mult_6/n790 ,
         \mul/mult_6/n789 , \mul/mult_6/n788 , \mul/mult_6/n787 ,
         \mul/mult_6/n786 , \mul/mult_6/n784 , \mul/mult_6/n783 ,
         \mul/mult_6/n782 , \mul/mult_6/n781 , \mul/mult_6/n780 ,
         \mul/mult_6/n779 , \mul/mult_6/n778 , \mul/mult_6/n777 ,
         \mul/mult_6/n776 , \mul/mult_6/n775 , \mul/mult_6/n774 ,
         \mul/mult_6/n773 , \mul/mult_6/n772 , \mul/mult_6/n771 ,
         \mul/mult_6/n770 , \mul/mult_6/n769 , \mul/mult_6/n768 ,
         \mul/mult_6/n767 , \mul/mult_6/n766 , \mul/mult_6/n765 ,
         \mul/mult_6/n764 , \mul/mult_6/n763 , \mul/mult_6/n762 ,
         \mul/mult_6/n761 , \mul/mult_6/n760 , \mul/mult_6/n759 ,
         \mul/mult_6/n731 , \mul/mult_6/n730 , \mul/mult_6/n729 ,
         \mul/mult_6/n728 , \mul/mult_6/n727 , \mul/mult_6/n726 ,
         \mul/mult_6/n725 , \mul/mult_6/n724 , \mul/mult_6/n723 ,
         \mul/mult_6/n722 , \mul/mult_6/n721 , \mul/mult_6/n720 ,
         \mul/mult_6/n719 , \mul/mult_6/n718 , \mul/mult_6/n717 ,
         \mul/mult_6/n716 , \mul/mult_6/n715 , \mul/mult_6/n714 ,
         \mul/mult_6/n713 , \mul/mult_6/n712 , \mul/mult_6/n708 ,
         \mul/mult_6/n707 , \mul/mult_6/n706 , \mul/mult_6/n705 ,
         \mul/mult_6/n704 , \mul/mult_6/n703 , \mul/mult_6/n702 ,
         \mul/mult_6/n701 , \mul/mult_6/n700 , \mul/mult_6/n699 ,
         \mul/mult_6/n698 , \mul/mult_6/n697 , \mul/mult_6/n696 ,
         \mul/mult_6/n695 , \mul/mult_6/n693 , \mul/mult_6/n692 ,
         \mul/mult_6/n691 , \mul/mult_6/n690 , \mul/mult_6/n689 ,
         \mul/mult_6/n688 , \mul/mult_6/n687 , \mul/mult_6/n686 ,
         \mul/mult_6/n685 , \mul/mult_6/n684 , \mul/mult_6/n683 ,
         \mul/mult_6/n682 , \mul/mult_6/n681 , \mul/mult_6/n680 ,
         \mul/mult_6/n679 , \mul/mult_6/n678 , \mul/mult_6/n677 ,
         \mul/mult_6/n676 , \mul/mult_6/n675 , \mul/mult_6/n674 ,
         \mul/mult_6/n673 , \mul/mult_6/n672 , \mul/mult_6/n671 ,
         \mul/mult_6/n670 , \mul/mult_6/n669 , \mul/mult_6/n668 ,
         \mul/mult_6/n667 , \mul/mult_6/n666 , \mul/mult_6/n665 ,
         \mul/mult_6/n664 , \mul/mult_6/n662 , \mul/mult_6/n661 ,
         \mul/mult_6/n660 , \mul/mult_6/n659 , \mul/mult_6/n658 ,
         \mul/mult_6/n655 , \mul/mult_6/n654 , \mul/mult_6/n653 ,
         \mul/mult_6/n652 , \mul/mult_6/n651 , \mul/mult_6/n650 ,
         \mul/mult_6/n649 , \mul/mult_6/n648 , \mul/mult_6/n646 ,
         \mul/mult_6/n645 , \mul/mult_6/n644 , \mul/mult_6/n643 ,
         \mul/mult_6/n640 , \mul/mult_6/n639 , \mul/mult_6/n638 ,
         \mul/mult_6/n637 , \mul/mult_6/n636 , \mul/mult_6/n635 ,
         \mul/mult_6/n634 , \mul/mult_6/n632 , \mul/mult_6/n631 ,
         \mul/mult_6/n630 , \mul/mult_6/n629 , \mul/mult_6/n628 ,
         \mul/mult_6/n627 , \mul/mult_6/n626 , \mul/mult_6/n625 ,
         \mul/mult_6/n624 , \mul/mult_6/n623 , \mul/mult_6/n622 ,
         \mul/mult_6/n621 , \mul/mult_6/n620 , \mul/mult_6/n619 ,
         \mul/mult_6/n617 , \mul/mult_6/n616 , \mul/mult_6/n615 ,
         \mul/mult_6/n614 , \mul/mult_6/n613 , \mul/mult_6/n612 ,
         \mul/mult_6/n611 , \mul/mult_6/n610 , \mul/mult_6/n609 ,
         \mul/mult_6/n608 , \mul/mult_6/n607 , \mul/mult_6/n605 ,
         \mul/mult_6/n604 , \mul/mult_6/n603 , \mul/mult_6/n602 ,
         \mul/mult_6/n601 , \mul/mult_6/n600 , \mul/mult_6/n599 ,
         \mul/mult_6/n598 , \mul/mult_6/n597 , \mul/mult_6/n596 ,
         \mul/mult_6/n595 , \mul/mult_6/n593 , \mul/mult_6/n592 ,
         \mul/mult_6/n591 , \mul/mult_6/n590 , \mul/mult_6/n589 ,
         \mul/mult_6/n588 , \mul/mult_6/n587 , \mul/mult_6/n585 ,
         \mul/mult_6/n583 , \mul/mult_6/n582 , \mul/mult_6/n581 ,
         \mul/mult_6/n580 , \mul/mult_6/n579 , \mul/mult_6/n576 ,
         \mul/mult_6/n575 , \mul/mult_6/n572 , \mul/mult_6/n571 ,
         \mul/mult_6/n570 , \mul/mult_6/n569 , \mul/mult_6/n568 ,
         \mul/mult_6/n567 , \mul/mult_6/n566 , \mul/mult_6/n565 ,
         \mul/mult_6/n564 , \mul/mult_6/n563 , \mul/mult_6/n562 ,
         \mul/mult_6/n561 , \mul/mult_6/n560 , \mul/mult_6/n559 ,
         \mul/mult_6/n558 , \mul/mult_6/n557 , \mul/mult_6/n556 ,
         \mul/mult_6/n555 , \mul/mult_6/n554 , \mul/mult_6/n553 ,
         \mul/mult_6/n552 , \mul/mult_6/n548 , \mul/mult_6/n547 ,
         \mul/mult_6/n544 , \mul/mult_6/n543 , \mul/mult_6/n540 ,
         \mul/mult_6/n539 , \mul/mult_6/n536 , \mul/mult_6/n535 ,
         \mul/mult_6/n532 , \mul/mult_6/n531 , \mul/mult_6/n528 ,
         \mul/mult_6/n524 , \mul/mult_6/n520 , \mul/mult_6/n495 ,
         \mul/mult_6/n494 , \mul/mult_6/n493 , \mul/mult_6/n492 ,
         \mul/mult_6/n491 , \mul/mult_6/n490 , \mul/mult_6/n489 ,
         \mul/mult_6/n488 , \mul/mult_6/n487 , \mul/mult_6/n486 ,
         \mul/mult_6/n485 , \mul/mult_6/n484 , \mul/mult_6/n483 ,
         \mul/mult_6/n482 , \mul/mult_6/n481 , \mul/mult_6/n480 ,
         \mul/mult_6/n479 , \mul/mult_6/n478 , \mul/mult_6/n477 ,
         \mul/mult_6/n476 , \mul/mult_6/n475 , \mul/mult_6/n474 ,
         \mul/mult_6/n473 , \mul/mult_6/n472 , \mul/mult_6/n471 ,
         \mul/mult_6/n470 , \mul/mult_6/n469 , \mul/mult_6/n468 ,
         \mul/mult_6/n467 , \mul/mult_6/n466 , \mul/mult_6/n465 ,
         \mul/mult_6/n464 , \mul/mult_6/n463 , \mul/mult_6/n462 ,
         \mul/mult_6/n461 , \mul/mult_6/n460 , \mul/mult_6/n459 ,
         \mul/mult_6/n458 , \mul/mult_6/n457 , \mul/mult_6/n456 ,
         \mul/mult_6/n455 , \mul/mult_6/n454 , \mul/mult_6/n453 ,
         \mul/mult_6/n452 , \mul/mult_6/n451 , \mul/mult_6/n450 ,
         \mul/mult_6/n449 , \mul/mult_6/n448 , \mul/mult_6/n447 ,
         \mul/mult_6/n446 , \mul/mult_6/n445 , \mul/mult_6/n444 ,
         \mul/mult_6/n443 , \mul/mult_6/n442 , \mul/mult_6/n441 ,
         \mul/mult_6/n440 , \mul/mult_6/n439 , \mul/mult_6/n438 ,
         \mul/mult_6/n437 , \mul/mult_6/n436 , \mul/mult_6/n435 ,
         \mul/mult_6/n434 , \mul/mult_6/n433 , \mul/mult_6/n432 ,
         \mul/mult_6/n431 , \mul/mult_6/n430 , \mul/mult_6/n429 ,
         \mul/mult_6/n428 , \mul/mult_6/n427 , \mul/mult_6/n426 ,
         \mul/mult_6/n425 , \mul/mult_6/n424 , \mul/mult_6/n423 ,
         \mul/mult_6/n422 , \mul/mult_6/n421 , \mul/mult_6/n420 ,
         \mul/mult_6/n419 , \mul/mult_6/n418 , \mul/mult_6/n417 ,
         \mul/mult_6/n416 , \mul/mult_6/n415 , \mul/mult_6/n414 ,
         \mul/mult_6/n413 , \mul/mult_6/n412 , \mul/mult_6/n411 ,
         \mul/mult_6/n410 , \mul/mult_6/n409 , \mul/mult_6/n408 ,
         \mul/mult_6/n407 , \mul/mult_6/n406 , \mul/mult_6/n405 ,
         \mul/mult_6/n404 , \mul/mult_6/n403 , \mul/mult_6/n402 ,
         \mul/mult_6/n401 , \mul/mult_6/n400 , \mul/mult_6/n399 ,
         \mul/mult_6/n398 , \mul/mult_6/n397 , \mul/mult_6/n396 ,
         \mul/mult_6/n395 , \mul/mult_6/n394 , \mul/mult_6/n393 ,
         \mul/mult_6/n392 , \mul/mult_6/n391 , \mul/mult_6/n390 ,
         \mul/mult_6/n389 , \mul/mult_6/n388 , \mul/mult_6/n387 ,
         \mul/mult_6/n386 , \mul/mult_6/n385 , \mul/mult_6/n384 ,
         \mul/mult_6/n383 , \mul/mult_6/n382 , \mul/mult_6/n381 ,
         \mul/mult_6/n380 , \mul/mult_6/n379 , \mul/mult_6/n378 ,
         \mul/mult_6/n377 , \mul/mult_6/n376 , \mul/mult_6/n375 ,
         \mul/mult_6/n374 , \mul/mult_6/n373 , \mul/mult_6/n372 ,
         \mul/mult_6/n371 , \mul/mult_6/n370 , \mul/mult_6/n369 ,
         \mul/mult_6/n368 , \mul/mult_6/n367 , \mul/mult_6/n366 ,
         \mul/mult_6/n365 , \mul/mult_6/n364 , \mul/mult_6/n363 ,
         \mul/mult_6/n362 , \mul/mult_6/n361 , \mul/mult_6/n360 ,
         \mul/mult_6/n359 , \mul/mult_6/n358 , \mul/mult_6/n357 ,
         \mul/mult_6/n356 , \mul/mult_6/n355 , \mul/mult_6/n354 ,
         \mul/mult_6/n353 , \mul/mult_6/n352 , \mul/mult_6/n351 ,
         \mul/mult_6/n350 , \mul/mult_6/n349 , \mul/mult_6/n348 ,
         \mul/mult_6/n347 , \mul/mult_6/n346 , \mul/mult_6/n345 ,
         \mul/mult_6/n344 , \mul/mult_6/n343 , \mul/mult_6/n342 ,
         \mul/mult_6/n341 , \mul/mult_6/n340 , \mul/mult_6/n339 ,
         \mul/mult_6/n338 , \mul/mult_6/n337 , \mul/mult_6/n336 ,
         \mul/mult_6/n335 , \mul/mult_6/n334 , \mul/mult_6/n333 ,
         \mul/mult_6/n332 , \mul/mult_6/n331 , \mul/mult_6/n330 ,
         \mul/mult_6/n329 , \mul/mult_6/n328 , \mul/mult_6/n327 ,
         \mul/mult_6/n326 , \mul/mult_6/n325 , \mul/mult_6/n324 ,
         \mul/mult_6/n323 , \mul/mult_6/n322 , \mul/mult_6/n321 ,
         \mul/mult_6/n320 , \mul/mult_6/n319 , \mul/mult_6/n318 ,
         \mul/mult_6/n317 , \mul/mult_6/n316 , \mul/mult_6/n315 ,
         \mul/mult_6/n314 , \mul/mult_6/n313 , \mul/mult_6/n312 ,
         \mul/mult_6/n311 , \mul/mult_6/n310 , \mul/mult_6/n309 ,
         \mul/mult_6/n308 , \mul/mult_6/n307 , \mul/mult_6/n306 ,
         \mul/mult_6/n305 , \mul/mult_6/n304 , \mul/mult_6/n303 ,
         \mul/mult_6/n302 , \mul/mult_6/n301 , \mul/mult_6/n300 ,
         \mul/mult_6/n299 , \mul/mult_6/n298 , \mul/mult_6/n297 ,
         \mul/mult_6/n296 , \mul/mult_6/n295 , \mul/mult_6/n294 ,
         \mul/mult_6/n293 , \mul/mult_6/n292 , \mul/mult_6/n291 ,
         \mul/mult_6/n290 , \mul/mult_6/n289 , \mul/mult_6/n287 ,
         \mul/mult_6/n286 , \mul/mult_6/n285 , \mul/mult_6/n284 ,
         \mul/mult_6/n283 , \mul/mult_6/n282 , \mul/mult_6/n281 ,
         \mul/mult_6/n280 , \mul/mult_6/n279 , \mul/mult_6/n277 ,
         \mul/mult_6/n276 , \mul/mult_6/n275 , \mul/mult_6/n274 ,
         \mul/mult_6/n273 , \mul/mult_6/n272 , \mul/mult_6/n271 ,
         \mul/mult_6/n270 , \mul/mult_6/n269 , \mul/mult_6/n268 ,
         \mul/mult_6/n267 , \mul/mult_6/n266 , \mul/mult_6/n265 ,
         \mul/mult_6/n264 , \mul/mult_6/n263 , \mul/mult_6/n262 ,
         \mul/mult_6/n261 , \mul/mult_6/n260 , \mul/mult_6/n258 ,
         \mul/mult_6/n257 , \mul/mult_6/n256 , \mul/mult_6/n255 ,
         \mul/mult_6/n254 , \mul/mult_6/n253 , \mul/mult_6/n252 ,
         \mul/mult_6/n251 , \mul/mult_6/n249 , \mul/mult_6/n248 ,
         \mul/mult_6/n247 , \mul/mult_6/n246 , \mul/mult_6/n245 ,
         \mul/mult_6/n244 , \mul/mult_6/n243 , \mul/mult_6/n242 ,
         \mul/mult_6/n241 , \mul/mult_6/n240 , \mul/mult_6/n239 ,
         \mul/mult_6/n238 , \mul/mult_6/n237 , \mul/mult_6/n236 ,
         \mul/mult_6/n235 , \mul/mult_6/n234 , \mul/mult_6/n232 ,
         \mul/mult_6/n231 , \mul/mult_6/n230 , \mul/mult_6/n229 ,
         \mul/mult_6/n228 , \mul/mult_6/n227 , \mul/mult_6/n225 ,
         \mul/mult_6/n224 , \mul/mult_6/n223 , \mul/mult_6/n222 ,
         \mul/mult_6/n221 , \mul/mult_6/n220 , \mul/mult_6/n219 ,
         \mul/mult_6/n218 , \mul/mult_6/n217 , \mul/mult_6/n216 ,
         \mul/mult_6/n215 , \mul/mult_6/n214 , \mul/mult_6/n212 ,
         \mul/mult_6/n211 , \mul/mult_6/n210 , \mul/mult_6/n209 ,
         \mul/mult_6/n208 , \mul/mult_6/n206 , \mul/mult_6/n205 ,
         \mul/mult_6/n204 , \mul/mult_6/n203 , \mul/mult_6/n202 ,
         \mul/mult_6/n201 , \mul/mult_6/n200 , \mul/mult_6/n199 ,
         \mul/mult_6/n198 , \mul/mult_6/n197 , \mul/mult_6/n195 ,
         \mul/mult_6/n194 , \mul/mult_6/n193 , \mul/mult_6/n191 ,
         \mul/mult_6/n190 , \mul/mult_6/n189 , \mul/mult_6/n188 ,
         \mul/mult_6/n187 , \mul/mult_6/n186 , \mul/mult_6/n184 ,
         \mul/mult_6/n183 , \mul/mult_6/n181 , \mul/mult_6/n180 ,
         \mul/mult_6/n176 , \mul/mult_6/n175 , \mul/mult_6/n173 ,
         \mul/mult_6/n172 , \mul/mult_6/n171 , \mul/mult_6/n170 ,
         \mul/mult_6/n169 , \mul/mult_6/n168 , \mul/mult_6/n167 ,
         \mul/mult_6/n166 , \mul/mult_6/n165 , \mul/mult_6/n164 ,
         \mul/mult_6/n163 , \mul/mult_6/n162 , \mul/mult_6/n161 ,
         \mul/mult_6/n160 , \mul/mult_6/n159 , \mul/mult_6/n158 ,
         \mul/mult_6/n157 , \mul/mult_6/n156 , \mul/mult_6/n155 ,
         \mul/mult_6/n154 , \mul/mult_6/n153 , \mul/mult_6/n152 ,
         \mul/mult_6/n151 , \mul/mult_6/n150 , \mul/mult_6/n149 ,
         \mul/mult_6/n148 , \mul/mult_6/n147 , \mul/mult_6/n146 ,
         \mul/mult_6/n145 , \mul/mult_6/n144 , \mul/mult_6/n143 ,
         \mul/mult_6/n142 , \mul/mult_6/n141 , \mul/mult_6/n140 ,
         \mul/mult_6/n139 , \mul/mult_6/n138 , \mul/mult_6/n137 ,
         \mul/mult_6/n136 , \mul/mult_6/n135 , \mul/mult_6/n134 ,
         \mul/mult_6/n133 , \mul/mult_6/n132 , \mul/mult_6/n131 ,
         \mul/mult_6/n130 , \mul/mult_6/n129 , \mul/mult_6/n128 ,
         \mul/mult_6/n127 , \mul/mult_6/n126 , \mul/mult_6/n125 ,
         \mul/mult_6/n78 , \mul/mult_6/n76 , \mul/mult_6/n74 ,
         \mul/mult_6/n72 , \mul/mult_6/n70 , \mul/mult_6/n68 ,
         \mul/mult_6/n64 , \mul/mult_6/n62 , \mul/mult_6/n60 ,
         \mul/mult_6/n58 , \mul/mult_6/n54 , \mul/mult_6/n52 ,
         \mul/mult_6/n50 , \mul/mult_6/n48 , \mul/mult_6/n42 ,
         \mul/mult_6/n40 , \mul/mult_6/n38 , \mul/mult_6/n32 ,
         \mul/mult_6/n30 , \mul/mult_6/n28 , \mul/mult_6/n22 ,
         \mul/mult_6/n20 , \mul/mult_6/n18 , \mul/mult_6/n12 , \mul/mult_6/n9 ,
         \mul/mult_6/n8 , \mul/mult_6/n2 , \sigadd/add_9/n295 ,
         \sigadd/add_9/n293 , \sigadd/add_9/n291 , \sigadd/add_9/n289 ,
         \sigadd/add_9/n287 , \sigadd/add_9/n285 , \sigadd/add_9/n283 ,
         \sigadd/add_9/n281 , \sigadd/add_9/n279 , \sigadd/add_9/n277 ,
         \sigadd/add_9/n275 , \sigadd/add_9/n273 , \sigadd/add_9/n271 ,
         \sigadd/add_9/n269 , \sigadd/add_9/n267 , \sigadd/add_9/n265 ,
         \sigadd/add_9/n263 , \sigadd/add_9/n261 , \sigadd/add_9/n259 ,
         \sigadd/add_9/n257 , \sigadd/add_9/n255 , \sigadd/add_9/n253 ,
         \sigadd/add_9/n251 , \sigadd/add_9/n249 , \sigadd/add_9/n246 ,
         \sigadd/add_9/n244 , \sigadd/add_9/n243 , \sigadd/add_9/n242 ,
         \sigadd/add_9/n241 , \sigadd/add_9/n239 , \sigadd/add_9/n237 ,
         \sigadd/add_9/n236 , \sigadd/add_9/n235 , \sigadd/add_9/n234 ,
         \sigadd/add_9/n233 , \sigadd/add_9/n231 , \sigadd/add_9/n229 ,
         \sigadd/add_9/n228 , \sigadd/add_9/n227 , \sigadd/add_9/n226 ,
         \sigadd/add_9/n225 , \sigadd/add_9/n223 , \sigadd/add_9/n221 ,
         \sigadd/add_9/n220 , \sigadd/add_9/n219 , \sigadd/add_9/n218 ,
         \sigadd/add_9/n217 , \sigadd/add_9/n215 , \sigadd/add_9/n213 ,
         \sigadd/add_9/n212 , \sigadd/add_9/n211 , \sigadd/add_9/n210 ,
         \sigadd/add_9/n209 , \sigadd/add_9/n207 , \sigadd/add_9/n205 ,
         \sigadd/add_9/n204 , \sigadd/add_9/n203 , \sigadd/add_9/n202 ,
         \sigadd/add_9/n201 , \sigadd/add_9/n199 , \sigadd/add_9/n197 ,
         \sigadd/add_9/n196 , \sigadd/add_9/n195 , \sigadd/add_9/n194 ,
         \sigadd/add_9/n193 , \sigadd/add_9/n191 , \sigadd/add_9/n189 ,
         \sigadd/add_9/n188 , \sigadd/add_9/n187 , \sigadd/add_9/n186 ,
         \sigadd/add_9/n185 , \sigadd/add_9/n183 , \sigadd/add_9/n181 ,
         \sigadd/add_9/n180 , \sigadd/add_9/n179 , \sigadd/add_9/n178 ,
         \sigadd/add_9/n177 , \sigadd/add_9/n175 , \sigadd/add_9/n173 ,
         \sigadd/add_9/n172 , \sigadd/add_9/n171 , \sigadd/add_9/n170 ,
         \sigadd/add_9/n169 , \sigadd/add_9/n167 , \sigadd/add_9/n165 ,
         \sigadd/add_9/n164 , \sigadd/add_9/n163 , \sigadd/add_9/n162 ,
         \sigadd/add_9/n161 , \sigadd/add_9/n159 , \sigadd/add_9/n157 ,
         \sigadd/add_9/n156 , \sigadd/add_9/n155 , \sigadd/add_9/n154 ,
         \sigadd/add_9/n153 , \sigadd/add_9/n151 , \sigadd/add_9/n149 ,
         \sigadd/add_9/n148 , \sigadd/add_9/n147 , \sigadd/add_9/n146 ,
         \sigadd/add_9/n145 , \sigadd/add_9/n143 , \sigadd/add_9/n141 ,
         \sigadd/add_9/n140 , \sigadd/add_9/n139 , \sigadd/add_9/n138 ,
         \sigadd/add_9/n137 , \sigadd/add_9/n135 , \sigadd/add_9/n133 ,
         \sigadd/add_9/n132 , \sigadd/add_9/n131 , \sigadd/add_9/n130 ,
         \sigadd/add_9/n129 , \sigadd/add_9/n127 , \sigadd/add_9/n125 ,
         \sigadd/add_9/n124 , \sigadd/add_9/n123 , \sigadd/add_9/n122 ,
         \sigadd/add_9/n121 , \sigadd/add_9/n119 , \sigadd/add_9/n117 ,
         \sigadd/add_9/n116 , \sigadd/add_9/n115 , \sigadd/add_9/n114 ,
         \sigadd/add_9/n113 , \sigadd/add_9/n111 , \sigadd/add_9/n109 ,
         \sigadd/add_9/n108 , \sigadd/add_9/n107 , \sigadd/add_9/n106 ,
         \sigadd/add_9/n105 , \sigadd/add_9/n103 , \sigadd/add_9/n101 ,
         \sigadd/add_9/n100 , \sigadd/add_9/n99 , \sigadd/add_9/n98 ,
         \sigadd/add_9/n97 , \sigadd/add_9/n95 , \sigadd/add_9/n93 ,
         \sigadd/add_9/n92 , \sigadd/add_9/n91 , \sigadd/add_9/n90 ,
         \sigadd/add_9/n89 , \sigadd/add_9/n87 , \sigadd/add_9/n85 ,
         \sigadd/add_9/n84 , \sigadd/add_9/n83 , \sigadd/add_9/n82 ,
         \sigadd/add_9/n81 , \sigadd/add_9/n79 , \sigadd/add_9/n77 ,
         \sigadd/add_9/n76 , \sigadd/add_9/n75 , \sigadd/add_9/n74 ,
         \sigadd/add_9/n73 , \sigadd/add_9/n71 , \sigadd/add_9/n69 ,
         \sigadd/add_9/n68 , \sigadd/add_9/n67 , \sigadd/add_9/n66 ,
         \sigadd/add_9/n65 , \sigadd/add_9/n63 , \sigadd/add_9/n61 ,
         \sigadd/add_9/n60 , \sigadd/add_9/n59 , \sigadd/add_9/n58 ,
         \sigadd/add_9/n57 , \sigadd/add_9/n55 , \sigadd/add_9/n53 ,
         \sigadd/add_9/n52 , \sigadd/add_9/n50 , \sigadd/add_9/n49 ,
         \sigadd/add_9/n48 , \sigadd/add_9/n47 , \sigadd/add_9/n46 ,
         \sigadd/add_9/n45 , \sigadd/add_9/n44 , \sigadd/add_9/n43 ,
         \sigadd/add_9/n42 , \sigadd/add_9/n41 , \sigadd/add_9/n40 ,
         \sigadd/add_9/n39 , \sigadd/add_9/n38 , \sigadd/add_9/n37 ,
         \sigadd/add_9/n36 , \sigadd/add_9/n35 , \sigadd/add_9/n34 ,
         \sigadd/add_9/n33 , \sigadd/add_9/n32 , \sigadd/add_9/n31 ,
         \sigadd/add_9/n30 , \sigadd/add_9/n29 , \sigadd/add_9/n28 ,
         \sigadd/add_9/n27 , \sigadd/add_9/n26 , \sigadd/add_9/n25 ,
         \sigadd/add_9/n24 , \sigadd/add_9/n23 , \sigadd/add_9/n22 ,
         \sigadd/add_9/n21 , \sigadd/add_9/n20 , \sigadd/add_9/n19 ,
         \sigadd/add_9/n18 , \sigadd/add_9/n17 , \sigadd/add_9/n16 ,
         \sigadd/add_9/n15 , \sigadd/add_9/n14 , \sigadd/add_9/n13 ,
         \sigadd/add_9/n12 , \sigadd/add_9/n11 , \sigadd/add_9/n10 ,
         \sigadd/add_9/n9 , \sigadd/add_9/n8 , \sigadd/add_9/n7 ,
         \sigadd/add_9/n6 , \sigadd/add_9/n5 , \sigadd/add_9/n4 ,
         \sigadd/add_9/n3 , \sigadd/add_9/n2 , \sigadd/add_9/n1 ,
         \sigadd/sub_add_11_b0/B[49] , \sigadd/sub_add_11_b0/n98 ,
         \sigadd/sub_add_11_b0/n97 , \sigadd/sub_add_11_b0/n96 ,
         \sigadd/sub_add_11_b0/n95 , \sigadd/sub_add_11_b0/n48 ,
         \sigadd/sub_add_11_b0/n47 , \sigadd/sub_add_11_b0/n46 ,
         \sigadd/sub_add_11_b0/n45 , \sigadd/sub_add_11_b0/n44 ,
         \sigadd/sub_add_11_b0/n43 , \sigadd/sub_add_11_b0/n42 ,
         \sigadd/sub_add_11_b0/n41 , \sigadd/sub_add_11_b0/n40 ,
         \sigadd/sub_add_11_b0/n39 , \sigadd/sub_add_11_b0/n38 ,
         \sigadd/sub_add_11_b0/n37 , \sigadd/sub_add_11_b0/n36 ,
         \sigadd/sub_add_11_b0/n35 , \sigadd/sub_add_11_b0/n34 ,
         \sigadd/sub_add_11_b0/n33 , \sigadd/sub_add_11_b0/n32 ,
         \sigadd/sub_add_11_b0/n31 , \sigadd/sub_add_11_b0/n30 ,
         \sigadd/sub_add_11_b0/n29 , \sigadd/sub_add_11_b0/n28 ,
         \sigadd/sub_add_11_b0/n27 , \sigadd/sub_add_11_b0/n26 ,
         \sigadd/sub_add_11_b0/n25 , \sigadd/sub_add_11_b0/n24 ,
         \sigadd/sub_add_11_b0/n23 , \sigadd/sub_add_11_b0/n22 ,
         \sigadd/sub_add_11_b0/n21 , \sigadd/sub_add_11_b0/n20 ,
         \sigadd/sub_add_11_b0/n19 , \sigadd/sub_add_11_b0/n18 ,
         \sigadd/sub_add_11_b0/n17 , \sigadd/sub_add_11_b0/n16 ,
         \sigadd/sub_add_11_b0/n15 , \sigadd/sub_add_11_b0/n14 ,
         \sigadd/sub_add_11_b0/n13 , \sigadd/sub_add_11_b0/n12 ,
         \sigadd/sub_add_11_b0/n11 , \sigadd/sub_add_11_b0/n10 ,
         \sigadd/sub_add_11_b0/n9 , \sigadd/sub_add_11_b0/n8 ,
         \sigadd/sub_add_11_b0/n7 , \sigadd/sub_add_11_b0/n6 ,
         \sigadd/sub_add_11_b0/n5 , \sigadd/sub_add_11_b0/n4 ,
         \sigadd/sub_add_11_b0/n3 , \sigadd/sub_add_11_b0/n2 ,
         \sigadd/sub_add_11_b0/n1 , \selc/r299/A[47] , \selc/r299/A[46] ,
         \selc/r299/A[45] , \selc/r299/A[44] , \selc/r299/A[43] ,
         \selc/r299/A[42] , \selc/r299/A[41] , \selc/r299/A[40] ,
         \selc/r299/A[39] , \selc/r299/A[38] , \selc/r299/A[37] ,
         \selc/r299/A[36] , \selc/r299/A[35] , \selc/r299/A[34] ,
         \selc/r299/A[33] , \selc/r299/A[32] , \selc/r299/A[31] ,
         \selc/r299/A[30] , \selc/r299/A[29] , \selc/r299/A[28] ,
         \selc/r299/A[27] , \selc/r299/A[26] , \selc/r299/A[25] ,
         \selc/r299/A[24] , \selc/r299/A[23] , \selc/r299/A[22] ,
         \selc/r299/A[21] , \selc/r299/A[20] , \selc/r299/A[19] ,
         \selc/r299/A[18] , \selc/r299/A[17] , \selc/r299/A[16] ,
         \selc/r299/A[15] , \selc/r299/A[14] , \selc/r299/A[13] ,
         \selc/r299/A[12] , \selc/r299/A[11] , \selc/r299/A[10] ,
         \selc/r299/A[9] , \selc/r299/A[8] , \selc/r299/A[7] ,
         \selc/r299/A[6] , \selc/r299/A[5] , \selc/r299/A[4] ,
         \selc/r299/A[3] , \selc/r299/A[2] , \selc/r299/A[1] , \selc/r299/n48 ,
         \selc/r299/n47 , \selc/r299/n46 , \selc/r299/n45 , \selc/r299/n44 ,
         \selc/r299/n43 , \selc/r299/n42 , \selc/r299/n41 , \selc/r299/n40 ,
         \selc/r299/n39 , \selc/r299/n38 , \selc/r299/n37 , \selc/r299/n36 ,
         \selc/r299/n35 , \selc/r299/n34 , \selc/r299/n33 , \selc/r299/n32 ,
         \selc/r299/n31 , \selc/r299/n30 , \selc/r299/n29 , \selc/r299/n28 ,
         \selc/r299/n27 , \selc/r299/n26 , \selc/r299/n25 , \selc/r299/n24 ,
         \selc/r299/n23 , \selc/r299/n22 , \selc/r299/n21 , \selc/r299/n20 ,
         \selc/r299/n19 , \selc/r299/n18 , \selc/r299/n17 , \selc/r299/n16 ,
         \selc/r299/n15 , \selc/r299/n14 , \selc/r299/n13 , \selc/r299/n12 ,
         \selc/r299/n11 , \selc/r299/n10 , \selc/r299/n9 , \selc/r299/n8 ,
         \selc/r299/n7 , \selc/r299/n6 , \selc/r299/n5 , \selc/r299/n4 ,
         \selc/r299/n3 , \selc/r299/n2 , \selc/r299/n1 , \sub/r301/n17 ,
         \sub/r301/n13 , \sub/r301/n7 , \sub/r301/n6 , \sub/r301/n5 ,
         \sub/r301/n4 , \sub/r301/n3 , \sub/r301/n2 , \sub/r301/n1 ,
         \sub/sub_17/n15 , \sub/sub_17/n14 , \sub/sub_17/n10 , \sub/sub_17/n7 ,
         \sub/sub_17/n6 , \sub/sub_17/n5 , \sub/sub_17/n4 , \sub/sub_17/n3 ,
         \sub/sub_17/n2 , \sub/sub_17/n1 ,
         \expadd/add_0_root_sub_0_root_sub_8/B[7] ,
         \expadd/add_0_root_sub_0_root_sub_8/B[0] ,
         \expadd/add_0_root_sub_0_root_sub_8/n11 ,
         \expadd/add_0_root_sub_0_root_sub_8/n9 ,
         \expadd/add_0_root_sub_0_root_sub_8/n8 ,
         \expadd/add_0_root_sub_0_root_sub_8/n7 ,
         \expadd/add_0_root_sub_0_root_sub_8/n6 ,
         \expadd/add_0_root_sub_0_root_sub_8/n5 ,
         \expadd/add_0_root_sub_0_root_sub_8/n4 ,
         \expadd/add_0_root_sub_0_root_sub_8/n3 ,
         \expadd/add_0_root_sub_0_root_sub_8/n2 ,
         \expadd/add_0_root_sub_0_root_sub_8/n1 , n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061;
  wire   [7:0] exp_A;
  wire   [7:0] exp_B;
  wire   [7:0] exp_C;
  wire   [24:0] sig_A;
  wire   [24:0] sig_B;
  wire   [49:0] sig_C;
  wire   [7:0] exp_P;
  wire   [49:0] sig_P;
  wire   [7:0] sub_out;
  wire   [7:0] mux_out;
  wire   [49:0] sel_P;
  wire   [49:0] sel_C;
  wire   [49:0] ali_P;
  wire   [49:0] ali_C;
  wire   [49:0] add_out;
  wire   [26:0] norm_out;
  wire   [5:0] zero_cnt;
  assign sign_A = A[31];
  assign sign_B = B[31];
  assign exp_A[7] = A[30];
  assign exp_A[6] = A[29];
  assign exp_A[5] = A[28];
  assign exp_A[4] = A[27];
  assign exp_A[3] = A[26];
  assign exp_A[2] = A[25];
  assign exp_A[1] = A[24];
  assign exp_A[0] = A[23];
  assign exp_B[7] = B[30];
  assign exp_B[6] = B[29];
  assign exp_B[5] = B[28];
  assign exp_B[4] = B[27];
  assign exp_B[3] = B[26];
  assign exp_B[2] = B[25];
  assign exp_B[1] = B[24];
  assign exp_B[0] = B[23];
  assign exp_C[7] = C[30];
  assign exp_C[6] = C[29];
  assign exp_C[5] = C[28];
  assign exp_C[4] = C[27];
  assign exp_C[3] = C[26];
  assign exp_C[2] = C[25];
  assign exp_C[1] = C[24];
  assign exp_C[0] = C[23];
  assign sig_A[22] = A[22];
  assign sig_A[21] = A[21];
  assign sig_A[20] = A[20];
  assign sig_A[19] = A[19];
  assign sig_A[18] = A[18];
  assign sig_A[17] = A[17];
  assign sig_A[16] = A[16];
  assign sig_A[15] = A[15];
  assign sig_A[14] = A[14];
  assign sig_A[13] = A[13];
  assign sig_A[12] = A[12];
  assign sig_A[11] = A[11];
  assign sig_A[10] = A[10];
  assign sig_A[9] = A[9];
  assign sig_A[8] = A[8];
  assign sig_A[7] = A[7];
  assign sig_A[6] = A[6];
  assign sig_A[5] = A[5];
  assign sig_A[4] = A[4];
  assign sig_A[3] = A[3];
  assign sig_A[2] = A[2];
  assign sig_A[1] = A[1];
  assign sig_A[0] = A[0];
  assign sig_B[22] = B[22];
  assign sig_B[21] = B[21];
  assign sig_B[20] = B[20];
  assign sig_B[19] = B[19];
  assign sig_B[18] = B[18];
  assign sig_B[17] = B[17];
  assign sig_B[16] = B[16];
  assign sig_B[15] = B[15];
  assign sig_B[14] = B[14];
  assign sig_B[13] = B[13];
  assign sig_B[12] = B[12];
  assign sig_B[11] = B[11];
  assign sig_B[10] = B[10];
  assign sig_B[9] = B[9];
  assign sig_B[8] = B[8];
  assign sig_B[7] = B[7];
  assign sig_B[6] = B[6];
  assign sig_B[5] = B[5];
  assign sig_B[4] = B[4];
  assign sig_B[3] = B[3];
  assign sig_B[2] = B[2];
  assign sig_B[1] = B[1];
  assign sig_B[0] = B[0];
  assign sig_C[45] = C[22];
  assign sig_C[44] = C[21];
  assign sig_C[43] = C[20];
  assign sig_C[42] = C[19];
  assign sig_C[41] = C[18];
  assign sig_C[40] = C[17];
  assign sig_C[39] = C[16];
  assign sig_C[38] = C[15];
  assign sig_C[37] = C[14];
  assign sig_C[36] = C[13];
  assign sig_C[35] = C[12];
  assign sig_C[34] = C[11];
  assign sig_C[33] = C[10];
  assign sig_C[32] = C[9];
  assign sig_C[31] = C[8];
  assign sig_C[30] = C[7];
  assign sig_C[29] = C[6];
  assign sig_C[28] = C[5];
  assign sig_C[27] = C[4];
  assign sig_C[26] = C[3];
  assign sig_C[25] = C[2];
  assign sig_C[24] = C[1];
  assign sig_C[23] = C[0];
  assign \two_en[1]  = C[31];

  MXI2X1 \align/sra_11/U742  ( .A(\align/sra_11/n478 ), .B(\align/sra_11/n606 ), .S0(sub_out[3]), .Y(\align/sra_11/n667 ) );
  MX2X1 \align/sra_11/U741  ( .A(sel_C[32]), .B(sel_C[33]), .S0(n507), .Y(
        \align/sra_11/n742 ) );
  MX2X1 \align/sra_11/U740  ( .A(sel_C[34]), .B(sel_C[35]), .S0(n507), .Y(
        \align/sra_11/n739 ) );
  MX2X1 \align/sra_11/U739  ( .A(sel_C[36]), .B(sel_C[37]), .S0(n507), .Y(
        \align/sra_11/n740 ) );
  MX2X1 \align/sra_11/U738  ( .A(sel_C[38]), .B(sel_C[39]), .S0(n507), .Y(
        \align/sra_11/n737 ) );
  MXI2X1 \align/sra_11/U737  ( .A(\align/sra_11/n722 ), .B(\align/sra_11/n719 ), .S0(n511), .Y(\align/sra_11/n607 ) );
  MX2X1 \align/sra_11/U736  ( .A(sel_C[40]), .B(sel_C[41]), .S0(n507), .Y(
        \align/sra_11/n738 ) );
  MX2X1 \align/sra_11/U735  ( .A(sel_C[42]), .B(sel_C[43]), .S0(n507), .Y(
        \align/sra_11/n734 ) );
  MX2X1 \align/sra_11/U734  ( .A(sel_C[44]), .B(sel_C[45]), .S0(n507), .Y(
        \align/sra_11/n735 ) );
  MX2X1 \align/sra_11/U733  ( .A(sel_C[46]), .B(\two_en[1] ), .S0(n507), .Y(
        \align/sra_11/n732 ) );
  MXI2X1 \align/sra_11/U732  ( .A(\align/sra_11/n720 ), .B(\align/sra_11/n716 ), .S0(n511), .Y(\align/sra_11/n604 ) );
  MX2X1 \align/sra_11/U731  ( .A(\two_en[1] ), .B(\two_en[1] ), .S0(n507), .Y(
        \align/sra_11/n733 ) );
  MXI2X1 \align/sra_11/U730  ( .A(\align/sra_11/n717 ), .B(n723), .S0(n511), 
        .Y(\align/sra_11/n605 ) );
  MXI2X1 \align/sra_11/U729  ( .A(\align/sra_11/n668 ), .B(\align/sra_11/n666 ), .S0(n719), .Y(\align/sra_11/n560 ) );
  MXI2X1 \align/sra_11/U725  ( .A(\align/sra_11/n653 ), .B(\align/sra_11/n650 ), .S0(sub_out[3]), .Y(\align/sra_11/n595 ) );
  MXI2X1 \align/sra_11/U723  ( .A(\align/sra_11/n651 ), .B(\two_en[1] ), .S0(
        sub_out[3]), .Y(\align/sra_11/n596 ) );
  MXI2X1 \align/sra_11/U722  ( .A(\align/sra_11/n731 ), .B(\align/sra_11/n528 ), .S0(n515), .Y(\align/sra_11/n730 ) );
  MXI2X1 \align/sra_11/U721  ( .A(n722), .B(\align/sra_11/n730 ), .S0(n510), 
        .Y(\align/N64 ) );
  MX2X1 \align/sra_11/U719  ( .A(sel_C[33]), .B(sel_C[34]), .S0(n507), .Y(
        \align/sra_11/n702 ) );
  MX2X1 \align/sra_11/U718  ( .A(sel_C[35]), .B(sel_C[36]), .S0(n507), .Y(
        \align/sra_11/n703 ) );
  MX2X1 \align/sra_11/U717  ( .A(sel_C[37]), .B(sel_C[38]), .S0(n507), .Y(
        \align/sra_11/n700 ) );
  MX2X1 \align/sra_11/U716  ( .A(sel_C[39]), .B(sel_C[40]), .S0(n507), .Y(
        \align/sra_11/n701 ) );
  MX2X1 \align/sra_11/U715  ( .A(sel_C[41]), .B(sel_C[42]), .S0(n507), .Y(
        \align/sra_11/n698 ) );
  MXI2X1 \align/sra_11/U714  ( .A(\align/sra_11/n676 ), .B(\align/sra_11/n673 ), .S0(n511), .Y(\align/sra_11/n644 ) );
  MX2X1 \align/sra_11/U712  ( .A(sel_C[43]), .B(sel_C[44]), .S0(n507), .Y(
        \align/sra_11/n699 ) );
  MX2X1 \align/sra_11/U711  ( .A(sel_C[45]), .B(sel_C[46]), .S0(n507), .Y(
        \align/sra_11/n695 ) );
  MX2X1 \align/sra_11/U710  ( .A(\two_en[1] ), .B(\two_en[1] ), .S0(n507), .Y(
        \align/sra_11/n696 ) );
  MXI2X1 \align/sra_11/U709  ( .A(\align/sra_11/n674 ), .B(\align/sra_11/n671 ), .S0(n511), .Y(\align/sra_11/n645 ) );
  MXI2X1 \align/sra_11/U708  ( .A(\align/sra_11/n728 ), .B(\align/sra_11/n526 ), .S0(n515), .Y(\align/sra_11/n727 ) );
  MXI2X1 \align/sra_11/U707  ( .A(n720), .B(\align/sra_11/n727 ), .S0(n510), 
        .Y(\align/N65 ) );
  MXI2X1 \align/sra_11/U705  ( .A(\align/sra_11/n631 ), .B(\align/sra_11/n628 ), .S0(n506), .Y(\align/sra_11/n587 ) );
  MXI2X1 \align/sra_11/U703  ( .A(\align/sra_11/n629 ), .B(\two_en[1] ), .S0(
        n506), .Y(\align/sra_11/n588 ) );
  MXI2X1 \align/sra_11/U702  ( .A(\align/sra_11/n715 ), .B(\align/sra_11/n524 ), .S0(n515), .Y(\align/sra_11/n714 ) );
  MXI2X1 \align/sra_11/U701  ( .A(n720), .B(\align/sra_11/n714 ), .S0(n510), 
        .Y(\align/N66 ) );
  MXI2X1 \align/sra_11/U698  ( .A(\align/sra_11/n659 ), .B(\align/sra_11/n656 ), .S0(n511), .Y(\align/sra_11/n622 ) );
  MXI2X1 \align/sra_11/U696  ( .A(\align/sra_11/n623 ), .B(\two_en[1] ), .S0(
        n506), .Y(\align/sra_11/n584 ) );
  MXI2X1 \align/sra_11/U695  ( .A(\align/sra_11/n694 ), .B(\align/sra_11/n522 ), .S0(n515), .Y(\align/sra_11/n693 ) );
  MXI2X1 \align/sra_11/U694  ( .A(n720), .B(\align/sra_11/n693 ), .S0(n510), 
        .Y(\align/N67 ) );
  MXI2X1 \align/sra_11/U692  ( .A(\align/sra_11/n619 ), .B(\align/sra_11/n616 ), .S0(n506), .Y(\align/sra_11/n567 ) );
  MXI2X1 \align/sra_11/U690  ( .A(\align/sra_11/n617 ), .B(\two_en[1] ), .S0(
        n506), .Y(\align/sra_11/n568 ) );
  MXI2X1 \align/sra_11/U689  ( .A(\align/sra_11/n682 ), .B(\align/sra_11/n520 ), .S0(n515), .Y(\align/sra_11/n681 ) );
  MXI2X1 \align/sra_11/U688  ( .A(n720), .B(\align/sra_11/n681 ), .S0(n510), 
        .Y(\align/N68 ) );
  MXI2X1 \align/sra_11/U686  ( .A(\align/sra_11/n613 ), .B(\align/sra_11/n610 ), .S0(n506), .Y(\align/sra_11/n563 ) );
  MXI2X1 \align/sra_11/U684  ( .A(\align/sra_11/n611 ), .B(\two_en[1] ), .S0(
        n506), .Y(\align/sra_11/n564 ) );
  MXI2X1 \align/sra_11/U683  ( .A(\align/sra_11/n670 ), .B(\align/sra_11/n518 ), .S0(n515), .Y(\align/sra_11/n669 ) );
  MXI2X1 \align/sra_11/U682  ( .A(n720), .B(\align/sra_11/n669 ), .S0(n510), 
        .Y(\align/N69 ) );
  MXI2X1 \align/sra_11/U681  ( .A(\align/sra_11/n665 ), .B(\align/sra_11/n516 ), .S0(n515), .Y(\align/sra_11/n664 ) );
  MXI2X1 \align/sra_11/U680  ( .A(n720), .B(\align/sra_11/n664 ), .S0(n510), 
        .Y(\align/N70 ) );
  MXI2X1 \align/sra_11/U679  ( .A(\align/sra_11/n471 ), .B(\align/sra_11/n600 ), .S0(n506), .Y(\align/sra_11/n636 ) );
  MXI2X1 \align/sra_11/U678  ( .A(\align/sra_11/n658 ), .B(\align/sra_11/n659 ), .S0(n511), .Y(\align/sra_11/n601 ) );
  MXI2X1 \align/sra_11/U677  ( .A(\align/sra_11/n656 ), .B(\align/sra_11/n657 ), .S0(n511), .Y(\align/sra_11/n599 ) );
  MXI2X1 \align/sra_11/U675  ( .A(n720), .B(\align/sra_11/n654 ), .S0(n510), 
        .Y(\align/N71 ) );
  MXI2X1 \align/sra_11/U674  ( .A(\align/sra_11/n652 ), .B(\align/sra_11/n653 ), .S0(n506), .Y(\align/sra_11/n573 ) );
  MXI2X1 \align/sra_11/U673  ( .A(\align/sra_11/n650 ), .B(\align/sra_11/n651 ), .S0(n506), .Y(\align/sra_11/n571 ) );
  MXI2X1 \align/sra_11/U671  ( .A(n720), .B(\align/sra_11/n648 ), .S0(n510), 
        .Y(\align/N72 ) );
  MXI2X1 \align/sra_11/U670  ( .A(\align/sra_11/n646 ), .B(\align/sra_11/n647 ), .S0(n506), .Y(\align/sra_11/n537 ) );
  MXI2X1 \align/sra_11/U669  ( .A(\align/sra_11/n644 ), .B(\align/sra_11/n645 ), .S0(n506), .Y(\align/sra_11/n554 ) );
  MXI2X1 \align/sra_11/U667  ( .A(n721), .B(\align/sra_11/n642 ), .S0(n510), 
        .Y(\align/N73 ) );
  MXI2X1 \align/sra_11/U666  ( .A(\align/sra_11/n634 ), .B(n723), .S0(
        sub_out[4]), .Y(\align/sra_11/n558 ) );
  MXI2X1 \align/sra_11/U665  ( .A(n720), .B(\align/sra_11/n632 ), .S0(n510), 
        .Y(\align/N55 ) );
  MXI2X1 \align/sra_11/U664  ( .A(\align/sra_11/n630 ), .B(\align/sra_11/n631 ), .S0(n506), .Y(\align/sra_11/n510 ) );
  MXI2X1 \align/sra_11/U663  ( .A(\align/sra_11/n628 ), .B(\align/sra_11/n629 ), .S0(n506), .Y(\align/sra_11/n552 ) );
  MXI2X1 \align/sra_11/U661  ( .A(n721), .B(\align/sra_11/n626 ), .S0(n510), 
        .Y(\align/N74 ) );
  MXI2X1 \align/sra_11/U660  ( .A(\align/sra_11/n624 ), .B(\align/sra_11/n625 ), .S0(n506), .Y(\align/sra_11/n501 ) );
  MXI2X1 \align/sra_11/U659  ( .A(\align/sra_11/n622 ), .B(\align/sra_11/n623 ), .S0(n506), .Y(\align/sra_11/n550 ) );
  MXI2X1 \align/sra_11/U657  ( .A(n720), .B(\align/sra_11/n620 ), .S0(n510), 
        .Y(\align/N75 ) );
  MXI2X1 \align/sra_11/U656  ( .A(\align/sra_11/n618 ), .B(\align/sra_11/n619 ), .S0(n506), .Y(\align/sra_11/n492 ) );
  MXI2X1 \align/sra_11/U655  ( .A(\align/sra_11/n616 ), .B(\align/sra_11/n617 ), .S0(n506), .Y(\align/sra_11/n548 ) );
  MXI2X1 \align/sra_11/U653  ( .A(n721), .B(\align/sra_11/n614 ), .S0(n510), 
        .Y(\align/N76 ) );
  MXI2X1 \align/sra_11/U652  ( .A(\align/sra_11/n612 ), .B(\align/sra_11/n613 ), .S0(n506), .Y(\align/sra_11/n483 ) );
  MXI2X1 \align/sra_11/U651  ( .A(\align/sra_11/n610 ), .B(\align/sra_11/n611 ), .S0(n506), .Y(\align/sra_11/n546 ) );
  MXI2X1 \align/sra_11/U649  ( .A(n721), .B(\align/sra_11/n608 ), .S0(n510), 
        .Y(\align/N77 ) );
  MXI2X1 \align/sra_11/U648  ( .A(n721), .B(\align/sra_11/n602 ), .S0(n510), 
        .Y(\align/N78 ) );
  MXI2X1 \align/sra_11/U646  ( .A(n721), .B(\align/sra_11/n597 ), .S0(n510), 
        .Y(\align/N79 ) );
  MXI2X1 \align/sra_11/U644  ( .A(n721), .B(\align/sra_11/n593 ), .S0(n510), 
        .Y(\align/N80 ) );
  MXI2X1 \align/sra_11/U642  ( .A(n722), .B(\align/sra_11/n589 ), .S0(n510), 
        .Y(\align/N81 ) );
  MXI2X1 \align/sra_11/U640  ( .A(n722), .B(\align/sra_11/n585 ), .S0(n510), 
        .Y(\align/N82 ) );
  MXI2X1 \align/sra_11/U638  ( .A(n722), .B(\align/sra_11/n581 ), .S0(n510), 
        .Y(\align/N83 ) );
  MXI2X1 \align/sra_11/U630  ( .A(n722), .B(\align/sra_11/n565 ), .S0(n510), 
        .Y(\align/N84 ) );
  MXI2X1 \align/sra_11/U628  ( .A(n722), .B(\align/sra_11/n561 ), .S0(n510), 
        .Y(\align/N85 ) );
  MXI2X1 \align/sra_11/U627  ( .A(n722), .B(\align/sra_11/n559 ), .S0(n510), 
        .Y(\align/N86 ) );
  MXI2X1 \align/sra_11/U625  ( .A(n722), .B(\align/sra_11/n557 ), .S0(n510), 
        .Y(\align/N87 ) );
  MXI2X1 \align/sra_11/U624  ( .A(n722), .B(\align/sra_11/n555 ), .S0(n510), 
        .Y(\align/N88 ) );
  MXI2X1 \align/sra_11/U623  ( .A(n722), .B(\align/sra_11/n553 ), .S0(n510), 
        .Y(\align/N89 ) );
  MXI2X1 \align/sra_11/U622  ( .A(n722), .B(\align/sra_11/n551 ), .S0(n510), 
        .Y(\align/N90 ) );
  MXI2X1 \align/sra_11/U621  ( .A(n721), .B(\align/sra_11/n549 ), .S0(n510), 
        .Y(\align/N91 ) );
  MXI2X1 \align/sra_11/U620  ( .A(n721), .B(\align/sra_11/n547 ), .S0(n510), 
        .Y(\align/N92 ) );
  MXI2X1 \align/sra_11/U619  ( .A(n721), .B(\align/sra_11/n545 ), .S0(n510), 
        .Y(\align/N93 ) );
  MXI2X1 \align/sra_11/U614  ( .A(n721), .B(\align/sra_11/n533 ), .S0(n510), 
        .Y(\align/N57 ) );
  MXI2X1 \align/sra_11/U613  ( .A(n721), .B(\align/sra_11/n531 ), .S0(n510), 
        .Y(\align/N94 ) );
  MXI2X1 \align/sra_11/U612  ( .A(n721), .B(\align/sra_11/n529 ), .S0(n510), 
        .Y(\align/N95 ) );
  MXI2X1 \align/sra_11/U611  ( .A(n722), .B(\align/sra_11/n527 ), .S0(n510), 
        .Y(\align/N96 ) );
  MXI2X1 \align/sra_11/U610  ( .A(n721), .B(\align/sra_11/n525 ), .S0(n510), 
        .Y(\align/N97 ) );
  MXI2X1 \align/sra_11/U609  ( .A(n721), .B(\align/sra_11/n523 ), .S0(n510), 
        .Y(\align/N98 ) );
  MXI2X1 \align/sra_11/U608  ( .A(n721), .B(\align/sra_11/n521 ), .S0(n510), 
        .Y(\align/N99 ) );
  MXI2X1 \align/sra_11/U607  ( .A(n723), .B(\align/sra_11/n519 ), .S0(n510), 
        .Y(\align/N100 ) );
  MXI2X1 \align/sra_11/U606  ( .A(n720), .B(\align/sra_11/n517 ), .S0(n510), 
        .Y(\align/N101 ) );
  MXI2X1 \align/sra_11/U605  ( .A(n723), .B(\align/sra_11/n515 ), .S0(n510), 
        .Y(\align/N102 ) );
  MXI2X1 \align/sra_11/U601  ( .A(\align/sra_11/n507 ), .B(\align/sra_11/n508 ), .S0(n515), .Y(\align/sra_11/n506 ) );
  MXI2X1 \align/sra_11/U600  ( .A(n722), .B(\align/sra_11/n506 ), .S0(n510), 
        .Y(\align/N58 ) );
  MXI2X1 \align/sra_11/U596  ( .A(\align/sra_11/n498 ), .B(\align/sra_11/n499 ), .S0(n515), .Y(\align/sra_11/n497 ) );
  MXI2X1 \align/sra_11/U595  ( .A(n722), .B(\align/sra_11/n497 ), .S0(n510), 
        .Y(\align/N59 ) );
  MXI2X1 \align/sra_11/U591  ( .A(\align/sra_11/n489 ), .B(\align/sra_11/n490 ), .S0(n515), .Y(\align/sra_11/n488 ) );
  MXI2X1 \align/sra_11/U590  ( .A(n721), .B(\align/sra_11/n488 ), .S0(n510), 
        .Y(\align/N60 ) );
  MXI2X1 \align/sra_11/U586  ( .A(\align/sra_11/n480 ), .B(\align/sra_11/n481 ), .S0(n515), .Y(\align/sra_11/n479 ) );
  MXI2X1 \align/sra_11/U585  ( .A(n721), .B(\align/sra_11/n479 ), .S0(n510), 
        .Y(\align/N61 ) );
  MXI2X1 \align/sra_11/U582  ( .A(\align/sra_11/n473 ), .B(\align/sra_11/n474 ), .S0(n515), .Y(\align/sra_11/n472 ) );
  MXI2X1 \align/sra_11/U581  ( .A(n720), .B(\align/sra_11/n472 ), .S0(n510), 
        .Y(\align/N62 ) );
  MXI2X1 \align/sra_11/U578  ( .A(\align/sra_11/n466 ), .B(\align/sra_11/n467 ), .S0(n515), .Y(\align/sra_11/n464 ) );
  MXI2X1 \align/sra_11/U577  ( .A(n722), .B(\align/sra_11/n464 ), .S0(n510), 
        .Y(\align/N63 ) );
  MX2X1 \align/sra_11/U405  ( .A(sel_C[24]), .B(sel_C[25]), .S0(n507), .Y(
        \align/sra_11/n746 ) );
  MXI2X1 \align/sra_11/U402  ( .A(\align/sra_11/n702 ), .B(\align/sra_11/n703 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n658 ) );
  MXI2X1 \align/sra_11/U401  ( .A(\align/sra_11/n733 ), .B(\two_en[1] ), .S0(
        \align/sra_11/SH[1] ), .Y(\align/sra_11/n717 ) );
  MXI2X1 \align/sra_11/U400  ( .A(\align/sra_11/n742 ), .B(\align/sra_11/n739 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n722 ) );
  MXI2X1 \align/sra_11/U399  ( .A(\align/sra_11/n738 ), .B(\align/sra_11/n734 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n720 ) );
  MXI2X1 \align/sra_11/U398  ( .A(\align/sra_11/n740 ), .B(\align/sra_11/n737 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n719 ) );
  MXI2X1 \align/sra_11/U397  ( .A(\align/sra_11/n735 ), .B(\align/sra_11/n732 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n716 ) );
  MXI2X1 \align/sra_11/U395  ( .A(\align/sra_11/n695 ), .B(\align/sra_11/n696 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n657 ) );
  MXI2X1 \align/sra_11/U394  ( .A(\align/sra_11/n698 ), .B(\align/sra_11/n699 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n656 ) );
  MXI2X1 \align/sra_11/U393  ( .A(\align/sra_11/n700 ), .B(\align/sra_11/n701 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n659 ) );
  MXI2X1 \align/sra_11/U392  ( .A(\align/sra_11/n706 ), .B(\align/sra_11/n707 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n660 ) );
  MXI2X1 \align/sra_11/U379  ( .A(\align/sra_11/n605 ), .B(\two_en[1] ), .S0(
        n506), .Y(\align/sra_11/n666 ) );
  MXI2X1 \align/sra_11/U378  ( .A(\align/sra_11/n554 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n535 ) );
  MXI2X1 \align/sra_11/U377  ( .A(\align/sra_11/n596 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n528 ) );
  MXI2X1 \align/sra_11/U376  ( .A(\align/sra_11/n588 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n524 ) );
  MXI2X1 \align/sra_11/U375  ( .A(\align/sra_11/n552 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n508 ) );
  MXI2X1 \align/sra_11/U374  ( .A(\align/sra_11/n607 ), .B(\align/sra_11/n604 ), .S0(n506), .Y(\align/sra_11/n668 ) );
  MXI2X1 \align/sra_11/U373  ( .A(\align/sra_11/n592 ), .B(n722), .S0(n719), 
        .Y(\align/sra_11/n526 ) );
  MXI2X1 \align/sra_11/U372  ( .A(\align/sra_11/n564 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n518 ) );
  MXI2X1 \align/sra_11/U371  ( .A(\align/sra_11/n530 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n467 ) );
  MXI2X1 \align/sra_11/U370  ( .A(\align/sra_11/n532 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n474 ) );
  MXI2X1 \align/sra_11/U369  ( .A(\align/sra_11/n546 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n481 ) );
  MXI2X1 \align/sra_11/U368  ( .A(\align/sra_11/n548 ), .B(n722), .S0(n719), 
        .Y(\align/sra_11/n490 ) );
  MXI2X1 \align/sra_11/U367  ( .A(\align/sra_11/n550 ), .B(n723), .S0(n719), 
        .Y(\align/sra_11/n499 ) );
  MXI2X1 \align/sra_11/U366  ( .A(\align/sra_11/n571 ), .B(n723), .S0(
        sub_out[4]), .Y(\align/sra_11/n556 ) );
  MXI2X1 \align/sra_11/U365  ( .A(\align/sra_11/n601 ), .B(\align/sra_11/n599 ), .S0(n506), .Y(\align/sra_11/n634 ) );
  AOI21X1 \mul/mult_6/U339  ( .A0(\mul/mult_6/n78 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n74 ), .Y(\mul/mult_6/n974 ) );
  OAI21X1 \mul/mult_6/U972  ( .A0(n544), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1355 ), .Y(\mul/mult_6/n1329 ) );
  XOR2X1 \sub/sub_17/U2  ( .A(\sub/sub_17/n10 ), .B(exp_C[7]), .Y(
        \sub/sub_17/n1 ) );
  XOR2X1 \sub/sub_17/U1  ( .A(\sub/sub_17/n2 ), .B(\sub/sub_17/n1 ), .Y(
        \sub/N21 ) );
  XOR2X1 \sub/r301/U1  ( .A(\sub/r301/n2 ), .B(\sub/r301/n1 ), .Y(\sub/N12 )
         );
  MXI2X1 \align/sra_10/U352  ( .A(sel_P[1]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n256 ) );
  MXI2X1 \align/sra_10/U351  ( .A(sel_P[2]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n257 ) );
  MXI2X1 \align/sra_10/U298  ( .A(\align/sra_10/n256 ), .B(\align/sra_10/n257 ), .S0(n507), .Y(\align/sra_10/n202 ) );
  MXI2X1 \align/sra_10/U350  ( .A(sel_P[3]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n258 ) );
  MXI2X1 \align/sra_10/U349  ( .A(sel_P[4]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n259 ) );
  MXI2X1 \align/sra_10/U296  ( .A(\align/sra_10/n258 ), .B(\align/sra_10/n259 ), .S0(n507), .Y(\align/sra_10/n204 ) );
  MXI2X1 \align/sra_10/U348  ( .A(sel_P[5]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n260 ) );
  MXI2X1 \align/sra_10/U347  ( .A(sel_P[6]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n261 ) );
  MXI2X1 \align/sra_10/U294  ( .A(\align/sra_10/n260 ), .B(\align/sra_10/n261 ), .S0(n507), .Y(\align/sra_10/n206 ) );
  MXI2X1 \align/sra_10/U346  ( .A(sel_P[7]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n262 ) );
  MXI2X1 \align/sra_10/U345  ( .A(sel_P[8]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n263 ) );
  MXI2X1 \align/sra_10/U292  ( .A(\align/sra_10/n262 ), .B(\align/sra_10/n263 ), .S0(n507), .Y(\align/sra_10/n208 ) );
  MXI2X1 \align/sra_10/U244  ( .A(\align/sra_10/n206 ), .B(\align/sra_10/n208 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n156 ) );
  MXI2X1 \align/sra_10/U198  ( .A(\align/sra_10/n152 ), .B(\align/sra_10/n156 ), .S0(n505), .Y(\align/sra_10/n102 ) );
  MXI2X1 \align/sra_10/U344  ( .A(sel_P[9]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n264 ) );
  MXI2X1 \align/sra_10/U343  ( .A(sel_P[10]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n265 ) );
  MXI2X1 \align/sra_10/U290  ( .A(\align/sra_10/n264 ), .B(\align/sra_10/n265 ), .S0(n507), .Y(\align/sra_10/n210 ) );
  MXI2X1 \align/sra_10/U342  ( .A(sel_P[11]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n266 ) );
  MXI2X1 \align/sra_10/U341  ( .A(sel_P[12]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n267 ) );
  MXI2X1 \align/sra_10/U288  ( .A(\align/sra_10/n266 ), .B(\align/sra_10/n267 ), .S0(n507), .Y(\align/sra_10/n212 ) );
  MXI2X1 \align/sra_10/U240  ( .A(\align/sra_10/n210 ), .B(\align/sra_10/n212 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n160 ) );
  MXI2X1 \align/sra_10/U340  ( .A(sel_P[13]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n268 ) );
  MXI2X1 \align/sra_10/U339  ( .A(sel_P[14]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n269 ) );
  MXI2X1 \align/sra_10/U286  ( .A(\align/sra_10/n268 ), .B(\align/sra_10/n269 ), .S0(n507), .Y(\align/sra_10/n214 ) );
  MXI2X1 \align/sra_10/U338  ( .A(sel_P[15]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n270 ) );
  MXI2X1 \align/sra_10/U337  ( .A(sel_P[16]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n271 ) );
  MXI2X1 \align/sra_10/U284  ( .A(\align/sra_10/n270 ), .B(\align/sra_10/n271 ), .S0(n507), .Y(\align/sra_10/n216 ) );
  MXI2X1 \align/sra_10/U236  ( .A(\align/sra_10/n214 ), .B(\align/sra_10/n216 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n164 ) );
  MXI2X1 \align/sra_10/U190  ( .A(\align/sra_10/n160 ), .B(\align/sra_10/n164 ), .S0(n505), .Y(\align/sra_10/n110 ) );
  MXI2X1 \align/sra_10/U148  ( .A(\align/sra_10/n102 ), .B(\align/sra_10/n110 ), .S0(n506), .Y(\align/sra_10/n52 ) );
  MXI2X1 \align/sra_10/U336  ( .A(sel_P[17]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n272 ) );
  MXI2X1 \align/sra_10/U335  ( .A(sel_P[18]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n273 ) );
  MXI2X1 \align/sra_10/U282  ( .A(\align/sra_10/n272 ), .B(\align/sra_10/n273 ), .S0(n507), .Y(\align/sra_10/n218 ) );
  MXI2X1 \align/sra_10/U334  ( .A(sel_P[19]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n274 ) );
  MXI2X1 \align/sra_10/U333  ( .A(sel_P[20]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n275 ) );
  MXI2X1 \align/sra_10/U280  ( .A(\align/sra_10/n274 ), .B(\align/sra_10/n275 ), .S0(n507), .Y(\align/sra_10/n220 ) );
  MXI2X1 \align/sra_10/U232  ( .A(\align/sra_10/n218 ), .B(\align/sra_10/n220 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n168 ) );
  MXI2X1 \align/sra_10/U332  ( .A(sel_P[21]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n276 ) );
  MXI2X1 \align/sra_10/U278  ( .A(\align/sra_10/n276 ), .B(\align/sra_10/n277 ), .S0(n507), .Y(\align/sra_10/n222 ) );
  MXI2X1 \align/sra_10/U330  ( .A(sel_P[23]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n278 ) );
  MXI2X1 \align/sra_10/U182  ( .A(\align/sra_10/n168 ), .B(\align/sra_10/n172 ), .S0(n505), .Y(\align/sra_10/n118 ) );
  MXI2X1 \align/sra_10/U328  ( .A(sel_P[25]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n280 ) );
  MXI2X1 \align/sra_10/U325  ( .A(sel_P[28]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n283 ) );
  MXI2X1 \align/sra_10/U132  ( .A(\align/sra_10/n118 ), .B(\align/sra_10/n126 ), .S0(n506), .Y(\align/sra_10/n68 ) );
  MX2X1 \align/sra_10/U48  ( .A(\align/sra_10/n2 ), .B(\align/sra_10/n18 ), 
        .S0(n719), .Y(\align/N5 ) );
  MX2X1 \align/sra_11/U521  ( .A(sel_C[23]), .B(sel_C[24]), .S0(n507), .Y(
        \align/sra_11/n709 ) );
  MX2X1 \align/sra_11/U527  ( .A(sel_C[25]), .B(sel_C[26]), .S0(n507), .Y(
        \align/sra_11/n706 ) );
  MX2X1 \align/sra_11/U525  ( .A(sel_C[27]), .B(sel_C[28]), .S0(n507), .Y(
        \align/sra_11/n707 ) );
  MX2X1 \align/sra_11/U528  ( .A(sel_C[29]), .B(sel_C[30]), .S0(n507), .Y(
        \align/sra_11/n704 ) );
  MX2X1 \align/sra_11/U526  ( .A(sel_C[31]), .B(sel_C[32]), .S0(n507), .Y(
        \align/sra_11/n705 ) );
  MXI2X1 \align/sra_11/U485  ( .A(\align/sra_11/n704 ), .B(\align/sra_11/n705 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n661 ) );
  MXI2X1 \align/sra_11/U450  ( .A(\align/sra_11/n660 ), .B(\align/sra_11/n661 ), .S0(n511), .Y(\align/sra_11/n600 ) );
  MXI2X1 \align/sra_10/U299  ( .A(\align/sra_10/n255 ), .B(\align/sra_10/n256 ), .S0(n507), .Y(\align/sra_10/n201 ) );
  MXI2X1 \align/sra_10/U297  ( .A(\align/sra_10/n257 ), .B(\align/sra_10/n258 ), .S0(n507), .Y(\align/sra_10/n203 ) );
  MXI2X1 \align/sra_10/U295  ( .A(\align/sra_10/n259 ), .B(\align/sra_10/n260 ), .S0(n507), .Y(\align/sra_10/n205 ) );
  MXI2X1 \align/sra_10/U293  ( .A(\align/sra_10/n261 ), .B(\align/sra_10/n262 ), .S0(n507), .Y(\align/sra_10/n207 ) );
  MXI2X1 \align/sra_10/U245  ( .A(\align/sra_10/n205 ), .B(\align/sra_10/n207 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n155 ) );
  MXI2X1 \align/sra_10/U291  ( .A(\align/sra_10/n263 ), .B(\align/sra_10/n264 ), .S0(n507), .Y(\align/sra_10/n209 ) );
  MXI2X1 \align/sra_10/U289  ( .A(\align/sra_10/n265 ), .B(\align/sra_10/n266 ), .S0(n507), .Y(\align/sra_10/n211 ) );
  MXI2X1 \align/sra_10/U241  ( .A(\align/sra_10/n209 ), .B(\align/sra_10/n211 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n159 ) );
  MXI2X1 \align/sra_10/U287  ( .A(\align/sra_10/n267 ), .B(\align/sra_10/n268 ), .S0(n507), .Y(\align/sra_10/n213 ) );
  MXI2X1 \align/sra_10/U285  ( .A(\align/sra_10/n269 ), .B(\align/sra_10/n270 ), .S0(n507), .Y(\align/sra_10/n215 ) );
  MXI2X1 \align/sra_10/U237  ( .A(\align/sra_10/n213 ), .B(\align/sra_10/n215 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n163 ) );
  MXI2X1 \align/sra_10/U191  ( .A(\align/sra_10/n159 ), .B(\align/sra_10/n163 ), .S0(n505), .Y(\align/sra_10/n109 ) );
  MXI2X1 \align/sra_10/U283  ( .A(\align/sra_10/n271 ), .B(\align/sra_10/n272 ), .S0(n507), .Y(\align/sra_10/n217 ) );
  MXI2X1 \align/sra_10/U281  ( .A(\align/sra_10/n273 ), .B(\align/sra_10/n274 ), .S0(n507), .Y(\align/sra_10/n219 ) );
  MXI2X1 \align/sra_10/U233  ( .A(\align/sra_10/n217 ), .B(\align/sra_10/n219 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n167 ) );
  MXI2X1 \align/sra_10/U279  ( .A(\align/sra_10/n275 ), .B(\align/sra_10/n276 ), .S0(n507), .Y(\align/sra_10/n221 ) );
  MXI2X1 \align/sra_10/U183  ( .A(\align/sra_10/n167 ), .B(\align/sra_10/n171 ), .S0(n505), .Y(\align/sra_10/n117 ) );
  MX2X1 \align/sra_11/U522  ( .A(sel_C[26]), .B(sel_C[27]), .S0(n507), .Y(
        \align/sra_11/n743 ) );
  MXI2X1 \align/sra_11/U483  ( .A(\align/sra_11/n746 ), .B(\align/sra_11/n743 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n724 ) );
  MX2X1 \align/sra_11/U524  ( .A(sel_C[28]), .B(sel_C[29]), .S0(n507), .Y(
        \align/sra_11/n744 ) );
  MX2X1 \align/sra_11/U523  ( .A(sel_C[30]), .B(sel_C[31]), .S0(n507), .Y(
        \align/sra_11/n741 ) );
  MXI2X1 \align/sra_11/U484  ( .A(\align/sra_11/n744 ), .B(\align/sra_11/n741 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n721 ) );
  MXI2X1 \align/sra_11/U449  ( .A(\align/sra_11/n724 ), .B(\align/sra_11/n721 ), .S0(n511), .Y(\align/sra_11/n606 ) );
  MXI2X1 \align/sra_10/U247  ( .A(\align/sra_10/n203 ), .B(\align/sra_10/n205 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n153 ) );
  MXI2X1 \align/sra_10/U243  ( .A(\align/sra_10/n207 ), .B(\align/sra_10/n209 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n157 ) );
  MXI2X1 \align/sra_10/U197  ( .A(\align/sra_10/n153 ), .B(\align/sra_10/n157 ), .S0(n505), .Y(\align/sra_10/n103 ) );
  MXI2X1 \align/sra_10/U239  ( .A(\align/sra_10/n211 ), .B(\align/sra_10/n213 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n161 ) );
  MXI2X1 \align/sra_10/U235  ( .A(\align/sra_10/n215 ), .B(\align/sra_10/n217 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n165 ) );
  MXI2X1 \align/sra_10/U189  ( .A(\align/sra_10/n161 ), .B(\align/sra_10/n165 ), .S0(n505), .Y(\align/sra_10/n111 ) );
  MXI2X1 \align/sra_10/U147  ( .A(\align/sra_10/n103 ), .B(\align/sra_10/n111 ), .S0(n506), .Y(\align/sra_10/n53 ) );
  MXI2X1 \align/sra_10/U231  ( .A(\align/sra_10/n219 ), .B(\align/sra_10/n221 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n169 ) );
  MXI2X1 \align/sra_10/U131  ( .A(\align/sra_10/n119 ), .B(\align/sra_10/n127 ), .S0(n506), .Y(\align/sra_10/n69 ) );
  MX2X1 \align/sra_10/U47  ( .A(\align/sra_10/n3 ), .B(\align/sra_10/n19 ), 
        .S0(n719), .Y(\align/N6 ) );
  MXI2X1 \align/sra_11/U492  ( .A(n653), .B(\align/sra_11/n746 ), .S0(
        \align/sra_11/SH[1] ), .Y(\align/sra_11/n689 ) );
  MXI2X1 \align/sra_11/U490  ( .A(\align/sra_11/n743 ), .B(\align/sra_11/n744 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n690 ) );
  MXI2X1 \align/sra_11/U491  ( .A(\align/sra_11/n741 ), .B(\align/sra_11/n742 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n687 ) );
  MXI2X1 \align/sra_11/U453  ( .A(\align/sra_11/n690 ), .B(\align/sra_11/n687 ), .S0(n511), .Y(\align/sra_11/n653 ) );
  MXI2X1 \align/sra_11/U488  ( .A(\align/sra_11/n739 ), .B(\align/sra_11/n740 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n688 ) );
  MXI2X1 \align/sra_11/U489  ( .A(\align/sra_11/n737 ), .B(\align/sra_11/n738 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n685 ) );
  MXI2X1 \align/sra_11/U452  ( .A(\align/sra_11/n688 ), .B(\align/sra_11/n685 ), .S0(n511), .Y(\align/sra_11/n650 ) );
  MXI2X1 \align/sra_11/U486  ( .A(\align/sra_11/n734 ), .B(\align/sra_11/n735 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n686 ) );
  MXI2X1 \align/sra_11/U487  ( .A(\align/sra_11/n732 ), .B(\align/sra_11/n733 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n683 ) );
  MXI2X1 \align/sra_11/U451  ( .A(\align/sra_11/n686 ), .B(\align/sra_11/n683 ), .S0(n511), .Y(\align/sra_11/n651 ) );
  XNOR2X1 \sigadd/add_9/U328  ( .A(\sigadd/add_9/n242 ), .B(\sigadd/add_9/n48 ), .Y(\sigadd/sig[2] ) );
  MXI2X1 \align/sra_10/U246  ( .A(\align/sra_10/n204 ), .B(\align/sra_10/n206 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n154 ) );
  MXI2X1 \align/sra_10/U242  ( .A(\align/sra_10/n208 ), .B(\align/sra_10/n210 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n158 ) );
  MXI2X1 \align/sra_10/U196  ( .A(\align/sra_10/n154 ), .B(\align/sra_10/n158 ), .S0(n505), .Y(\align/sra_10/n104 ) );
  MXI2X1 \align/sra_10/U238  ( .A(\align/sra_10/n212 ), .B(\align/sra_10/n214 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n162 ) );
  MXI2X1 \align/sra_10/U234  ( .A(\align/sra_10/n216 ), .B(\align/sra_10/n218 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n166 ) );
  MXI2X1 \align/sra_10/U188  ( .A(\align/sra_10/n162 ), .B(\align/sra_10/n166 ), .S0(n505), .Y(\align/sra_10/n112 ) );
  MXI2X1 \align/sra_10/U146  ( .A(\align/sra_10/n104 ), .B(\align/sra_10/n112 ), .S0(n506), .Y(\align/sra_10/n54 ) );
  MXI2X1 \align/sra_10/U230  ( .A(\align/sra_10/n220 ), .B(\align/sra_10/n222 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n170 ) );
  MXI2X1 \align/sra_10/U130  ( .A(\align/sra_10/n120 ), .B(\align/sra_10/n128 ), .S0(n506), .Y(\align/sra_10/n70 ) );
  MX2X1 \align/sra_10/U46  ( .A(\align/sra_10/n4 ), .B(\align/sra_10/n20 ), 
        .S0(n718), .Y(\align/N7 ) );
  MXI2X1 \align/sra_11/U494  ( .A(\align/sra_11/n709 ), .B(\align/sra_11/n706 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n677 ) );
  MXI2X1 \align/sra_11/U498  ( .A(\align/sra_11/n707 ), .B(\align/sra_11/n704 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n678 ) );
  MXI2X1 \align/sra_11/U499  ( .A(\align/sra_11/n705 ), .B(\align/sra_11/n702 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n675 ) );
  MXI2X1 \align/sra_11/U455  ( .A(\align/sra_11/n678 ), .B(\align/sra_11/n675 ), .S0(n511), .Y(\align/sra_11/n647 ) );
  MXI2X1 \align/sra_11/U493  ( .A(\align/sra_11/n703 ), .B(\align/sra_11/n700 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n676 ) );
  MXI2X1 \align/sra_11/U496  ( .A(\align/sra_11/n701 ), .B(\align/sra_11/n698 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n673 ) );
  MXI2X1 \align/sra_11/U495  ( .A(\align/sra_11/n699 ), .B(\align/sra_11/n695 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_11/n674 ) );
  MXI2X1 \align/sra_11/U497  ( .A(\align/sra_11/n696 ), .B(\two_en[1] ), .S0(
        \align/sra_11/SH[1] ), .Y(\align/sra_11/n671 ) );
  MXI2X1 \align/sra_10/U195  ( .A(\align/sra_10/n155 ), .B(\align/sra_10/n159 ), .S0(n505), .Y(\align/sra_10/n105 ) );
  MXI2X1 \align/sra_10/U187  ( .A(\align/sra_10/n163 ), .B(\align/sra_10/n167 ), .S0(n505), .Y(\align/sra_10/n113 ) );
  MXI2X1 \align/sra_10/U145  ( .A(\align/sra_10/n105 ), .B(\align/sra_10/n113 ), .S0(n506), .Y(\align/sra_10/n55 ) );
  MXI2X1 \align/sra_10/U95  ( .A(\align/sra_10/n55 ), .B(\align/sra_10/n87 ), 
        .S0(n717), .Y(\align/sra_10/n5 ) );
  MX2X1 \align/sra_10/U45  ( .A(\align/sra_10/n5 ), .B(\align/sra_10/n21 ), 
        .S0(n718), .Y(\align/N8 ) );
  MXI2X1 \align/sra_11/U460  ( .A(\align/sra_11/n723 ), .B(\align/sra_11/n724 ), .S0(n511), .Y(\align/sra_11/n630 ) );
  MXI2X1 \align/sra_11/U459  ( .A(\align/sra_11/n721 ), .B(\align/sra_11/n722 ), .S0(n511), .Y(\align/sra_11/n631 ) );
  MXI2X1 \align/sra_11/U458  ( .A(\align/sra_11/n719 ), .B(\align/sra_11/n720 ), .S0(n511), .Y(\align/sra_11/n628 ) );
  MXI2X1 \align/sra_11/U457  ( .A(\align/sra_11/n716 ), .B(\align/sra_11/n717 ), .S0(n511), .Y(\align/sra_11/n629 ) );
  MXI2X1 \align/sra_10/U194  ( .A(\align/sra_10/n156 ), .B(\align/sra_10/n160 ), .S0(n505), .Y(\align/sra_10/n106 ) );
  MXI2X1 \align/sra_10/U186  ( .A(\align/sra_10/n164 ), .B(\align/sra_10/n168 ), .S0(n505), .Y(\align/sra_10/n114 ) );
  MXI2X1 \align/sra_10/U144  ( .A(\align/sra_10/n106 ), .B(\align/sra_10/n114 ), .S0(n506), .Y(\align/sra_10/n56 ) );
  MXI2X1 \align/sra_10/U94  ( .A(\align/sra_10/n56 ), .B(\align/sra_10/n88 ), 
        .S0(n717), .Y(\align/sra_10/n6 ) );
  MX2X1 \align/sra_10/U44  ( .A(\align/sra_10/n6 ), .B(\align/sra_10/n22 ), 
        .S0(n718), .Y(\align/N9 ) );
  MXI2X1 \align/sra_11/U463  ( .A(\align/sra_11/n663 ), .B(\align/sra_11/n660 ), .S0(n511), .Y(\align/sra_11/n624 ) );
  MXI2X1 \align/sra_11/U462  ( .A(\align/sra_11/n661 ), .B(\align/sra_11/n658 ), .S0(n511), .Y(\align/sra_11/n625 ) );
  MXI2X1 \align/sra_11/U461  ( .A(\align/sra_11/n657 ), .B(n720), .S0(n511), 
        .Y(\align/sra_11/n623 ) );
  MXI2X1 \align/sra_10/U193  ( .A(\align/sra_10/n157 ), .B(\align/sra_10/n161 ), .S0(n505), .Y(\align/sra_10/n107 ) );
  MXI2X1 \align/sra_10/U185  ( .A(\align/sra_10/n165 ), .B(\align/sra_10/n169 ), .S0(n505), .Y(\align/sra_10/n115 ) );
  MXI2X1 \align/sra_10/U143  ( .A(\align/sra_10/n107 ), .B(\align/sra_10/n115 ), .S0(n506), .Y(\align/sra_10/n57 ) );
  MXI2X1 \align/sra_10/U93  ( .A(\align/sra_10/n57 ), .B(\align/sra_10/n89 ), 
        .S0(n717), .Y(\align/sra_10/n7 ) );
  MXI2X1 \align/sra_11/U468  ( .A(\align/sra_11/n689 ), .B(\align/sra_11/n690 ), .S0(n511), .Y(\align/sra_11/n618 ) );
  MXI2X1 \align/sra_11/U467  ( .A(\align/sra_11/n687 ), .B(\align/sra_11/n688 ), .S0(n511), .Y(\align/sra_11/n619 ) );
  MXI2X1 \align/sra_11/U466  ( .A(\align/sra_11/n685 ), .B(\align/sra_11/n686 ), .S0(n511), .Y(\align/sra_11/n616 ) );
  MXI2X1 \align/sra_11/U465  ( .A(\align/sra_11/n683 ), .B(n720), .S0(n511), 
        .Y(\align/sra_11/n617 ) );
  MXI2X1 \align/sra_10/U192  ( .A(\align/sra_10/n158 ), .B(\align/sra_10/n162 ), .S0(n505), .Y(\align/sra_10/n108 ) );
  MXI2X1 \align/sra_10/U184  ( .A(\align/sra_10/n166 ), .B(\align/sra_10/n170 ), .S0(n505), .Y(\align/sra_10/n116 ) );
  MXI2X1 \align/sra_10/U142  ( .A(\align/sra_10/n108 ), .B(\align/sra_10/n116 ), .S0(n506), .Y(\align/sra_10/n58 ) );
  MXI2X1 \align/sra_10/U92  ( .A(\align/sra_10/n58 ), .B(\align/sra_10/n90 ), 
        .S0(n515), .Y(\align/sra_10/n8 ) );
  MXI2X1 \align/sra_11/U472  ( .A(\align/sra_11/n677 ), .B(\align/sra_11/n678 ), .S0(n511), .Y(\align/sra_11/n612 ) );
  MXI2X1 \align/sra_11/U471  ( .A(\align/sra_11/n675 ), .B(\align/sra_11/n676 ), .S0(n511), .Y(\align/sra_11/n613 ) );
  MXI2X1 \align/sra_11/U469  ( .A(\align/sra_11/n673 ), .B(\align/sra_11/n674 ), .S0(n511), .Y(\align/sra_11/n610 ) );
  MXI2X1 \align/sra_11/U470  ( .A(\align/sra_11/n671 ), .B(n720), .S0(n511), 
        .Y(\align/sra_11/n611 ) );
  MXI2X1 \align/sra_10/U141  ( .A(\align/sra_10/n109 ), .B(\align/sra_10/n117 ), .S0(n506), .Y(\align/sra_10/n59 ) );
  MXI2X1 \align/sra_10/U91  ( .A(\align/sra_10/n59 ), .B(\align/sra_10/n91 ), 
        .S0(n515), .Y(\align/sra_10/n9 ) );
  MXI2X1 \align/sra_11/U407  ( .A(\align/sra_11/n606 ), .B(\align/sra_11/n607 ), .S0(sub_out[3]), .Y(\align/sra_11/n476 ) );
  MXI2X1 \align/sra_11/U406  ( .A(\align/sra_11/n604 ), .B(\align/sra_11/n605 ), .S0(sub_out[3]), .Y(\align/sra_11/n532 ) );
  MXI2X1 \align/sra_10/U140  ( .A(\align/sra_10/n110 ), .B(\align/sra_10/n118 ), .S0(n506), .Y(\align/sra_10/n60 ) );
  MXI2X1 \align/sra_10/U90  ( .A(\align/sra_10/n60 ), .B(\align/sra_10/n92 ), 
        .S0(n515), .Y(\align/sra_10/n10 ) );
  MXI2X1 \align/sra_11/U409  ( .A(\align/sra_11/n600 ), .B(\align/sra_11/n601 ), .S0(sub_out[3]), .Y(\align/sra_11/n469 ) );
  MXI2X1 \align/sra_11/U408  ( .A(\align/sra_11/n599 ), .B(\two_en[1] ), .S0(
        sub_out[3]), .Y(\align/sra_11/n530 ) );
  MXI2X1 \align/sra_10/U139  ( .A(\align/sra_10/n111 ), .B(\align/sra_10/n119 ), .S0(n506), .Y(\align/sra_10/n61 ) );
  MXI2X1 \align/sra_10/U89  ( .A(\align/sra_10/n61 ), .B(\align/sra_10/n93 ), 
        .S0(n515), .Y(\align/sra_10/n11 ) );
  MXI2X1 \align/sra_10/U138  ( .A(\align/sra_10/n112 ), .B(\align/sra_10/n120 ), .S0(n506), .Y(\align/sra_10/n62 ) );
  MXI2X1 \align/sra_10/U88  ( .A(\align/sra_10/n62 ), .B(\align/sra_10/n94 ), 
        .S0(n515), .Y(\align/sra_10/n12 ) );
  MXI2X1 \align/sra_11/U411  ( .A(\align/sra_11/n647 ), .B(\align/sra_11/n644 ), .S0(sub_out[3]), .Y(\align/sra_11/n591 ) );
  MXI2X1 \align/sra_11/U410  ( .A(\align/sra_11/n645 ), .B(\two_en[1] ), .S0(
        sub_out[3]), .Y(\align/sra_11/n592 ) );
  MXI2X1 \align/sra_10/U137  ( .A(\align/sra_10/n113 ), .B(\align/sra_10/n121 ), .S0(n506), .Y(\align/sra_10/n63 ) );
  MXI2X1 \align/sra_10/U87  ( .A(\align/sra_10/n63 ), .B(\align/sra_10/n95 ), 
        .S0(n515), .Y(\align/sra_10/n13 ) );
  MXI2X1 \align/sra_10/U136  ( .A(\align/sra_10/n114 ), .B(\align/sra_10/n122 ), .S0(n506), .Y(\align/sra_10/n64 ) );
  MXI2X1 \align/sra_10/U86  ( .A(\align/sra_10/n64 ), .B(\align/sra_10/n96 ), 
        .S0(sub_out[5]), .Y(\align/sra_10/n14 ) );
  MXI2X1 \align/sra_11/U413  ( .A(\align/sra_11/n625 ), .B(\align/sra_11/n622 ), .S0(sub_out[3]), .Y(\align/sra_11/n583 ) );
  MXI2X1 \align/sra_11/U412  ( .A(\align/sra_11/n584 ), .B(n720), .S0(n718), 
        .Y(\align/sra_11/n522 ) );
  MXI2X1 \align/sra_10/U135  ( .A(\align/sra_10/n115 ), .B(\align/sra_10/n123 ), .S0(n506), .Y(\align/sra_10/n65 ) );
  MXI2X1 \align/sra_10/U85  ( .A(\align/sra_10/n65 ), .B(\align/sra_10/n97 ), 
        .S0(n515), .Y(\align/sra_10/n15 ) );
  MXI2X1 \align/sra_11/U414  ( .A(\align/sra_11/n568 ), .B(n720), .S0(n718), 
        .Y(\align/sra_11/n520 ) );
  MXI2X1 \align/sra_10/U134  ( .A(\align/sra_10/n116 ), .B(\align/sra_10/n124 ), .S0(n506), .Y(\align/sra_10/n66 ) );
  MXI2X1 \align/sra_10/U84  ( .A(\align/sra_10/n66 ), .B(\align/sra_10/n98 ), 
        .S0(n717), .Y(\align/sra_10/n16 ) );
  MXI2X1 \align/sra_11/U416  ( .A(\align/sra_11/n667 ), .B(\align/sra_11/n668 ), .S0(n719), .Y(\align/sra_11/n665 ) );
  MXI2X1 \align/sra_11/U415  ( .A(\align/sra_11/n666 ), .B(n720), .S0(n718), 
        .Y(\align/sra_11/n516 ) );
  MXI2X1 \align/sra_11/U417  ( .A(\align/sra_11/n636 ), .B(\align/sra_11/n634 ), .S0(n719), .Y(\align/sra_11/n655 ) );
  MXI2X1 \align/sra_11/U418  ( .A(\align/sra_11/n573 ), .B(\align/sra_11/n571 ), .S0(n719), .Y(\align/sra_11/n649 ) );
  MXI2X1 \align/sra_11/U419  ( .A(\align/sra_11/n537 ), .B(\align/sra_11/n554 ), .S0(n718), .Y(\align/sra_11/n643 ) );
  MXI2X1 \align/sra_11/U420  ( .A(\align/sra_11/n510 ), .B(\align/sra_11/n552 ), .S0(n718), .Y(\align/sra_11/n627 ) );
  MXI2X1 \align/sra_11/U421  ( .A(\align/sra_11/n501 ), .B(\align/sra_11/n550 ), .S0(n718), .Y(\align/sra_11/n621 ) );
  MXI2X1 \align/sra_11/U422  ( .A(\align/sra_11/n492 ), .B(\align/sra_11/n548 ), .S0(n718), .Y(\align/sra_11/n615 ) );
  MXI2X1 \align/sra_11/U423  ( .A(\align/sra_11/n483 ), .B(\align/sra_11/n546 ), .S0(n718), .Y(\align/sra_11/n609 ) );
  MXI2X1 \align/sra_11/U425  ( .A(\align/sra_11/n476 ), .B(\align/sra_11/n532 ), .S0(n718), .Y(\align/sra_11/n603 ) );
  MXI2X1 \align/sra_11/U426  ( .A(\align/sra_11/n469 ), .B(\align/sra_11/n530 ), .S0(n718), .Y(\align/sra_11/n598 ) );
  MXI2X1 \align/sra_11/U427  ( .A(\align/sra_11/n595 ), .B(\align/sra_11/n596 ), .S0(n718), .Y(\align/sra_11/n594 ) );
  MXI2X1 \align/sra_11/U433  ( .A(\align/sra_11/n560 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n559 ) );
  MXI2X1 \align/sra_10/U50  ( .A(\align/sra_10/n100 ), .B(n508), .S0(n515), 
        .Y(\align/sra_10/n50 ) );
  MXI2X1 \align/sra_11/U435  ( .A(\align/sra_11/n535 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n553 ) );
  MXI2X1 \align/sra_11/U436  ( .A(\align/sra_11/n508 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n551 ) );
  MXI2X1 \align/sra_11/U437  ( .A(\align/sra_11/n499 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n549 ) );
  MXI2X1 \align/sra_11/U438  ( .A(\align/sra_11/n490 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n547 ) );
  MXI2X1 \align/sra_11/U439  ( .A(\align/sra_11/n481 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n545 ) );
  MXI2X1 \align/sra_11/U440  ( .A(\align/sra_11/n474 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n531 ) );
  XNOR2X1 \sigadd/add_9/U314  ( .A(\sigadd/add_9/n234 ), .B(\sigadd/add_9/n46 ), .Y(\sigadd/sig[4] ) );
  XOR2X1 \sigadd/add_9/U322  ( .A(\sigadd/add_9/n237 ), .B(\sigadd/add_9/n47 ), 
        .Y(\sigadd/sig[3] ) );
  MXI2X1 \normal/srl_15/U207  ( .A(\normal/srl_15/n236 ), .B(
        \normal/srl_15/n238 ), .S0(n715), .Y(\normal/srl_15/n186 ) );
  MXI2X1 \normal/srl_15/U199  ( .A(\normal/srl_15/n244 ), .B(
        \normal/srl_15/n246 ), .S0(n514), .Y(\normal/srl_15/n194 ) );
  MXI2X1 \normal/srl_15/U107  ( .A(\normal/srl_15/n136 ), .B(
        \normal/srl_15/n144 ), .S0(n513), .Y(\normal/srl_15/n86 ) );
  MXI2X1 \normal/srl_15/U203  ( .A(\normal/srl_15/n240 ), .B(
        \normal/srl_15/n242 ), .S0(n514), .Y(\normal/srl_15/n190 ) );
  MXI2X1 \normal/srl_15/U103  ( .A(\normal/srl_15/n140 ), .B(
        \normal/srl_15/n148 ), .S0(n513), .Y(\normal/srl_15/n90 ) );
  MXI2X1 \normal/srl_15/U57  ( .A(\normal/srl_15/n86 ), .B(\normal/srl_15/n90 ), .S0(n512), .Y(\normal/srl_15/n38 ) );
  MXI2X1 \normal/srl_15/U206  ( .A(\normal/srl_15/n237 ), .B(
        \normal/srl_15/n239 ), .S0(n715), .Y(\normal/srl_15/n187 ) );
  MXI2X1 \normal/srl_15/U198  ( .A(\normal/srl_15/n245 ), .B(
        \normal/srl_15/n247 ), .S0(n514), .Y(\normal/srl_15/n195 ) );
  MXI2X1 \normal/srl_15/U106  ( .A(\normal/srl_15/n137 ), .B(
        \normal/srl_15/n145 ), .S0(n513), .Y(\normal/srl_15/n87 ) );
  MXI2X1 \normal/srl_15/U202  ( .A(\normal/srl_15/n241 ), .B(
        \normal/srl_15/n243 ), .S0(n514), .Y(\normal/srl_15/n191 ) );
  MXI2X1 \normal/srl_15/U56  ( .A(\normal/srl_15/n87 ), .B(\normal/srl_15/n91 ), .S0(n512), .Y(\normal/srl_15/n39 ) );
  MXI2X1 \normal/sll_15/U244  ( .A(add_out[37]), .B(\normal/srl_15/A[21] ), 
        .S0(n703), .Y(\normal/sll_15/n226 ) );
  MXI2X1 \normal/sll_15/U246  ( .A(add_out[35]), .B(add_out[19]), .S0(n703), 
        .Y(\normal/sll_15/n224 ) );
  MXI2X1 \normal/sll_15/U197  ( .A(\normal/sll_15/n226 ), .B(
        \normal/sll_15/n224 ), .S0(n514), .Y(\normal/sll_15/n179 ) );
  MXI2X1 \normal/sll_15/U229  ( .A(\normal/sll_15/n194 ), .B(
        \normal/sll_15/n192 ), .S0(n514), .Y(\normal/sll_15/n147 ) );
  MXI2X1 \normal/sll_15/U150  ( .A(\normal/sll_15/n179 ), .B(
        \normal/sll_15/n147 ), .S0(n504), .Y(\normal/sll_15/n132 ) );
  MXI2X1 \normal/sll_15/U252  ( .A(\normal/srl_15/A[29] ), .B(add_out[13]), 
        .S0(n703), .Y(\normal/sll_15/n218 ) );
  MXI2X1 \normal/sll_15/U254  ( .A(\normal/srl_15/A[27] ), .B(
        \normal/srl_15/A[11] ), .S0(n703), .Y(\normal/sll_15/n216 ) );
  MXI2X1 \normal/sll_15/U103  ( .A(\normal/sll_15/n132 ), .B(
        \normal/sll_15/n124 ), .S0(n513), .Y(\normal/sll_15/n85 ) );
  MXI2X1 \normal/sll_15/U248  ( .A(add_out[33]), .B(add_out[17]), .S0(n703), 
        .Y(\normal/sll_15/n222 ) );
  MXI2X1 \normal/sll_15/U250  ( .A(add_out[31]), .B(add_out[15]), .S0(n703), 
        .Y(\normal/sll_15/n220 ) );
  MXI2X1 \normal/sll_15/U201  ( .A(\normal/sll_15/n222 ), .B(
        \normal/sll_15/n220 ), .S0(n715), .Y(\normal/sll_15/n175 ) );
  MXI2X1 \normal/sll_15/U154  ( .A(\normal/sll_15/n175 ), .B(
        \normal/sll_15/n143 ), .S0(n504), .Y(\normal/sll_15/n128 ) );
  MXI2X1 \normal/sll_15/U256  ( .A(\normal/srl_15/A[25] ), .B(
        \normal/srl_15/A[9] ), .S0(n703), .Y(\normal/sll_15/n214 ) );
  MXI2X1 \normal/sll_15/U258  ( .A(add_out[23]), .B(add_out[7]), .S0(n703), 
        .Y(\normal/sll_15/n212 ) );
  MXI2X1 \normal/sll_15/U209  ( .A(\normal/sll_15/n214 ), .B(
        \normal/sll_15/n212 ), .S0(n514), .Y(\normal/sll_15/n167 ) );
  MXI2X1 \normal/sll_15/U107  ( .A(\normal/sll_15/n128 ), .B(
        \normal/sll_15/n120 ), .S0(n513), .Y(\normal/sll_15/n81 ) );
  MXI2X1 \normal/sll_15/U56  ( .A(\normal/sll_15/n85 ), .B(\normal/sll_15/n81 ), .S0(n704), .Y(\normal/sll_15/n38 ) );
  MXI2X1 \normal/sll_15/U245  ( .A(\normal/srl_15/A[36] ), .B(add_out[20]), 
        .S0(n703), .Y(\normal/sll_15/n225 ) );
  MXI2X1 \normal/sll_15/U247  ( .A(add_out[34]), .B(add_out[18]), .S0(n703), 
        .Y(\normal/sll_15/n223 ) );
  MXI2X1 \normal/sll_15/U198  ( .A(\normal/sll_15/n225 ), .B(
        \normal/sll_15/n223 ), .S0(n514), .Y(\normal/sll_15/n178 ) );
  MXI2X1 \normal/sll_15/U230  ( .A(\normal/sll_15/n193 ), .B(
        \normal/sll_15/n191 ), .S0(n715), .Y(\normal/sll_15/n146 ) );
  MXI2X1 \normal/sll_15/U151  ( .A(\normal/sll_15/n178 ), .B(
        \normal/sll_15/n146 ), .S0(n504), .Y(\normal/sll_15/n131 ) );
  MXI2X1 \normal/sll_15/U253  ( .A(add_out[28]), .B(\normal/srl_15/A[12] ), 
        .S0(n703), .Y(\normal/sll_15/n217 ) );
  MXI2X1 \normal/sll_15/U255  ( .A(add_out[26]), .B(\normal/srl_15/A[10] ), 
        .S0(n703), .Y(\normal/sll_15/n215 ) );
  MXI2X1 \normal/sll_15/U206  ( .A(\normal/sll_15/n217 ), .B(
        \normal/sll_15/n215 ), .S0(n514), .Y(\normal/sll_15/n170 ) );
  MXI2X1 \normal/sll_15/U104  ( .A(\normal/sll_15/n131 ), .B(
        \normal/sll_15/n123 ), .S0(n513), .Y(\normal/sll_15/n84 ) );
  MXI2X1 \normal/sll_15/U249  ( .A(\normal/srl_15/A[32] ), .B(add_out[16]), 
        .S0(n703), .Y(\normal/sll_15/n221 ) );
  MXI2X1 \normal/sll_15/U251  ( .A(add_out[30]), .B(add_out[14]), .S0(n703), 
        .Y(\normal/sll_15/n219 ) );
  MXI2X1 \normal/sll_15/U202  ( .A(\normal/sll_15/n221 ), .B(
        \normal/sll_15/n219 ), .S0(n715), .Y(\normal/sll_15/n174 ) );
  MXI2X1 \normal/sll_15/U155  ( .A(\normal/sll_15/n174 ), .B(
        \normal/sll_15/n142 ), .S0(n504), .Y(\normal/sll_15/n127 ) );
  MXI2X1 \normal/sll_15/U257  ( .A(add_out[24]), .B(\normal/srl_15/A[8] ), 
        .S0(n703), .Y(\normal/sll_15/n213 ) );
  MXI2X1 \normal/sll_15/U259  ( .A(\normal/srl_15/A[22] ), .B(
        \normal/srl_15/A[6] ), .S0(n703), .Y(\normal/sll_15/n211 ) );
  MXI2X1 \normal/sll_15/U108  ( .A(\normal/sll_15/n127 ), .B(
        \normal/sll_15/n119 ), .S0(n513), .Y(\normal/sll_15/n80 ) );
  MXI2X1 \normal/sll_15/U57  ( .A(\normal/sll_15/n84 ), .B(\normal/sll_15/n80 ), .S0(n704), .Y(\normal/sll_15/n37 ) );
  MXI2X1 \normal/srl_15/U208  ( .A(\normal/srl_15/n235 ), .B(
        \normal/srl_15/n237 ), .S0(n715), .Y(\normal/srl_15/n185 ) );
  MXI2X1 \normal/srl_15/U200  ( .A(\normal/srl_15/n243 ), .B(
        \normal/srl_15/n245 ), .S0(n514), .Y(\normal/srl_15/n193 ) );
  MXI2X1 \normal/srl_15/U108  ( .A(\normal/srl_15/n135 ), .B(
        \normal/srl_15/n143 ), .S0(n513), .Y(\normal/srl_15/n85 ) );
  MXI2X1 \normal/srl_15/U204  ( .A(\normal/srl_15/n239 ), .B(
        \normal/srl_15/n241 ), .S0(n514), .Y(\normal/srl_15/n189 ) );
  MXI2X1 \normal/srl_15/U104  ( .A(\normal/srl_15/n139 ), .B(
        \normal/srl_15/n147 ), .S0(n513), .Y(\normal/srl_15/n89 ) );
  MXI2X1 \normal/srl_15/U58  ( .A(\normal/srl_15/n85 ), .B(\normal/srl_15/n89 ), .S0(n512), .Y(\normal/srl_15/n37 ) );
  MXI2X1 \normal/sll_15/U199  ( .A(\normal/sll_15/n224 ), .B(
        \normal/sll_15/n222 ), .S0(n514), .Y(\normal/sll_15/n177 ) );
  MXI2X1 \normal/sll_15/U231  ( .A(\normal/sll_15/n192 ), .B(
        \normal/sll_15/n190 ), .S0(n715), .Y(\normal/sll_15/n145 ) );
  MXI2X1 \normal/sll_15/U152  ( .A(\normal/sll_15/n177 ), .B(
        \normal/sll_15/n145 ), .S0(n504), .Y(\normal/sll_15/n130 ) );
  MXI2X1 \normal/sll_15/U207  ( .A(\normal/sll_15/n216 ), .B(
        \normal/sll_15/n214 ), .S0(n715), .Y(\normal/sll_15/n169 ) );
  MXI2X1 \normal/sll_15/U105  ( .A(\normal/sll_15/n130 ), .B(
        \normal/sll_15/n122 ), .S0(n513), .Y(\normal/sll_15/n83 ) );
  MXI2X1 \normal/sll_15/U203  ( .A(\normal/sll_15/n220 ), .B(
        \normal/sll_15/n218 ), .S0(n514), .Y(\normal/sll_15/n173 ) );
  MXI2X1 \normal/sll_15/U260  ( .A(\normal/srl_15/A[21] ), .B(add_out[5]), 
        .S0(n703), .Y(\normal/sll_15/n210 ) );
  MXI2X1 \normal/sll_15/U109  ( .A(\normal/sll_15/n126 ), .B(
        \normal/sll_15/n118 ), .S0(n513), .Y(\normal/sll_15/n79 ) );
  MXI2X1 \normal/srl_15/U205  ( .A(\normal/srl_15/n238 ), .B(
        \normal/srl_15/n240 ), .S0(n514), .Y(\normal/srl_15/n188 ) );
  MXI2X1 \normal/srl_15/U197  ( .A(\normal/srl_15/n246 ), .B(
        \normal/srl_15/n248 ), .S0(n514), .Y(\normal/srl_15/n196 ) );
  MXI2X1 \normal/srl_15/U105  ( .A(\normal/srl_15/n138 ), .B(
        \normal/srl_15/n146 ), .S0(n513), .Y(\normal/srl_15/n88 ) );
  MXI2X1 \normal/srl_15/U201  ( .A(\normal/srl_15/n242 ), .B(
        \normal/srl_15/n244 ), .S0(n514), .Y(\normal/srl_15/n192 ) );
  MXI2X1 \normal/srl_15/U55  ( .A(\normal/srl_15/n88 ), .B(\normal/srl_15/n92 ), .S0(n704), .Y(\normal/srl_15/n40 ) );
  MXI2X1 \normal/sll_15/U243  ( .A(add_out[38]), .B(\normal/srl_15/A[22] ), 
        .S0(n703), .Y(\normal/sll_15/n227 ) );
  MXI2X1 \normal/sll_15/U196  ( .A(\normal/sll_15/n227 ), .B(
        \normal/sll_15/n225 ), .S0(n514), .Y(\normal/sll_15/n180 ) );
  MXI2X1 \normal/sll_15/U228  ( .A(\normal/sll_15/n195 ), .B(
        \normal/sll_15/n193 ), .S0(n715), .Y(\normal/sll_15/n148 ) );
  MXI2X1 \normal/sll_15/U149  ( .A(\normal/sll_15/n180 ), .B(
        \normal/sll_15/n148 ), .S0(n504), .Y(\normal/sll_15/n133 ) );
  MXI2X1 \normal/sll_15/U102  ( .A(\normal/sll_15/n133 ), .B(
        \normal/sll_15/n125 ), .S0(n513), .Y(\normal/sll_15/n86 ) );
  MXI2X1 \normal/sll_15/U200  ( .A(\normal/sll_15/n223 ), .B(
        \normal/sll_15/n221 ), .S0(n514), .Y(\normal/sll_15/n176 ) );
  MXI2X1 \normal/sll_15/U232  ( .A(\normal/sll_15/n191 ), .B(
        \normal/sll_15/n189 ), .S0(n715), .Y(\normal/sll_15/n144 ) );
  MXI2X1 \normal/sll_15/U208  ( .A(\normal/sll_15/n215 ), .B(
        \normal/sll_15/n213 ), .S0(n715), .Y(\normal/sll_15/n168 ) );
  MXI2X1 \normal/sll_15/U106  ( .A(\normal/sll_15/n129 ), .B(
        \normal/sll_15/n121 ), .S0(n513), .Y(\normal/sll_15/n82 ) );
  MXI2X1 \normal/sll_15/U55  ( .A(\normal/sll_15/n86 ), .B(\normal/sll_15/n82 ), .S0(n704), .Y(\normal/sll_15/n39 ) );
  MXI2X1 \normal/srl_15/U54  ( .A(\normal/srl_15/n89 ), .B(\normal/srl_15/n93 ), .S0(n704), .Y(\normal/srl_15/n41 ) );
  MXI2X1 \normal/sll_15/U242  ( .A(add_out[39]), .B(add_out[23]), .S0(n703), 
        .Y(\normal/sll_15/n228 ) );
  MXI2X1 \normal/sll_15/U195  ( .A(\normal/sll_15/n228 ), .B(
        \normal/sll_15/n226 ), .S0(n514), .Y(\normal/sll_15/n181 ) );
  MXI2X1 \normal/sll_15/U227  ( .A(\normal/sll_15/n196 ), .B(
        \normal/sll_15/n194 ), .S0(n514), .Y(\normal/sll_15/n149 ) );
  MXI2X1 \normal/sll_15/U148  ( .A(\normal/sll_15/n181 ), .B(
        \normal/sll_15/n149 ), .S0(n504), .Y(\normal/sll_15/n134 ) );
  MXI2X1 \normal/sll_15/U101  ( .A(\normal/sll_15/n134 ), .B(
        \normal/sll_15/n126 ), .S0(n513), .Y(\normal/sll_15/n87 ) );
  MXI2X1 \normal/srl_15/U209  ( .A(\normal/srl_15/n234 ), .B(
        \normal/srl_15/n236 ), .S0(n715), .Y(\normal/srl_15/n184 ) );
  MXI2X1 \normal/srl_15/U109  ( .A(\normal/srl_15/n134 ), .B(
        \normal/srl_15/n142 ), .S0(n513), .Y(\normal/srl_15/n84 ) );
  MXI2X1 \normal/srl_15/U59  ( .A(\normal/srl_15/n84 ), .B(\normal/srl_15/n88 ), .S0(n512), .Y(\normal/srl_15/n36 ) );
  MXI2X1 \normal/sll_15/U261  ( .A(add_out[20]), .B(\normal/srl_15/A[4] ), 
        .S0(n714), .Y(\normal/sll_15/n209 ) );
  MXI2X1 \normal/sll_15/U110  ( .A(\normal/sll_15/n125 ), .B(
        \normal/sll_15/n117 ), .S0(n513), .Y(\normal/sll_15/n78 ) );
  MXI2X1 \normal/srl_15/U210  ( .A(\normal/srl_15/n233 ), .B(
        \normal/srl_15/n235 ), .S0(n715), .Y(\normal/srl_15/n183 ) );
  MXI2X1 \normal/srl_15/U110  ( .A(\normal/srl_15/n133 ), .B(
        \normal/srl_15/n141 ), .S0(n513), .Y(\normal/srl_15/n83 ) );
  MXI2X1 \normal/srl_15/U60  ( .A(\normal/srl_15/n83 ), .B(\normal/srl_15/n87 ), .S0(n512), .Y(\normal/srl_15/n35 ) );
  MXI2X1 \normal/sll_15/U262  ( .A(add_out[19]), .B(add_out[3]), .S0(n714), 
        .Y(\normal/sll_15/n208 ) );
  MXI2X1 \normal/sll_15/U111  ( .A(\normal/sll_15/n124 ), .B(
        \normal/sll_15/n116 ), .S0(n513), .Y(\normal/sll_15/n77 ) );
  MXI2X1 \normal/sll_15/U60  ( .A(\normal/sll_15/n81 ), .B(\normal/sll_15/n77 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n34 ) );
  MXI2X1 \normal/srl_15/U262  ( .A(\normal/srl_15/A[32] ), .B(add_out[48]), 
        .S0(n703), .Y(\normal/srl_15/n231 ) );
  MXI2X1 \normal/srl_15/U212  ( .A(\normal/srl_15/n231 ), .B(
        \normal/srl_15/n233 ), .S0(n715), .Y(\normal/srl_15/n181 ) );
  MXI2X1 \normal/srl_15/U112  ( .A(\normal/srl_15/n131 ), .B(
        \normal/srl_15/n139 ), .S0(n513), .Y(\normal/srl_15/n81 ) );
  MXI2X1 \normal/srl_15/U62  ( .A(\normal/srl_15/n81 ), .B(\normal/srl_15/n85 ), .S0(n512), .Y(\normal/srl_15/n33 ) );
  MXI2X1 \normal/srl_15/U261  ( .A(add_out[33]), .B(add_out[49]), .S0(n703), 
        .Y(\normal/srl_15/n232 ) );
  MXI2X1 \normal/srl_15/U211  ( .A(\normal/srl_15/n232 ), .B(
        \normal/srl_15/n234 ), .S0(n715), .Y(\normal/srl_15/n182 ) );
  MXI2X1 \normal/srl_15/U111  ( .A(\normal/srl_15/n132 ), .B(
        \normal/srl_15/n140 ), .S0(n513), .Y(\normal/srl_15/n82 ) );
  MXI2X1 \normal/srl_15/U61  ( .A(\normal/srl_15/n82 ), .B(\normal/srl_15/n86 ), .S0(n512), .Y(\normal/srl_15/n34 ) );
  MXI2X1 \normal/sll_15/U263  ( .A(add_out[18]), .B(add_out[2]), .S0(n714), 
        .Y(\normal/sll_15/n207 ) );
  MXI2X1 \normal/sll_15/U112  ( .A(\normal/sll_15/n123 ), .B(
        \normal/sll_15/n115 ), .S0(n513), .Y(\normal/sll_15/n76 ) );
  MXI2X1 \normal/sll_15/U61  ( .A(\normal/sll_15/n80 ), .B(\normal/sll_15/n76 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n33 ) );
  MXI2X1 \normal/sll_15/U264  ( .A(add_out[17]), .B(\normal/srl_15/A[1] ), 
        .S0(n714), .Y(\normal/sll_15/n206 ) );
  MXI2X1 \normal/sll_15/U113  ( .A(\normal/sll_15/n122 ), .B(
        \normal/sll_15/n114 ), .S0(n513), .Y(\normal/sll_15/n75 ) );
  MXI2X1 \normal/sll_15/U62  ( .A(\normal/sll_15/n79 ), .B(\normal/sll_15/n75 ), .S0(n704), .Y(\normal/sll_15/n32 ) );
  MXI2X1 \normal/srl_15/U264  ( .A(add_out[30]), .B(add_out[46]), .S0(n703), 
        .Y(\normal/srl_15/n229 ) );
  MXI2X1 \normal/srl_15/U114  ( .A(\normal/srl_15/n129 ), .B(
        \normal/srl_15/n137 ), .S0(n513), .Y(\normal/srl_15/n79 ) );
  MXI2X1 \normal/srl_15/U64  ( .A(\normal/srl_15/n79 ), .B(\normal/srl_15/n83 ), .S0(n512), .Y(\normal/srl_15/n31 ) );
  MXI2X1 \normal/srl_15/U263  ( .A(add_out[31]), .B(add_out[47]), .S0(n703), 
        .Y(\normal/srl_15/n230 ) );
  MXI2X1 \normal/srl_15/U113  ( .A(\normal/srl_15/n130 ), .B(
        \normal/srl_15/n138 ), .S0(n513), .Y(\normal/srl_15/n80 ) );
  MXI2X1 \normal/srl_15/U63  ( .A(\normal/srl_15/n80 ), .B(\normal/srl_15/n84 ), .S0(n512), .Y(\normal/srl_15/n32 ) );
  MXI2X1 \normal/srl_15/U17  ( .A(\normal/srl_15/n31 ), .B(\normal/srl_15/n32 ), .S0(n503), .Y(\normal/N32 ) );
  MXI2X1 \normal/sll_15/U265  ( .A(add_out[16]), .B(\sigadd/sig[0] ), .S0(n714), .Y(\normal/sll_15/n205 ) );
  MXI2X1 \normal/sll_15/U114  ( .A(\normal/sll_15/n121 ), .B(
        \normal/sll_15/n113 ), .S0(n513), .Y(\normal/sll_15/n74 ) );
  MXI2X1 \normal/sll_15/U63  ( .A(\normal/sll_15/n78 ), .B(\normal/sll_15/n74 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n31 ) );
  MXI2X1 \normal/sll_15/U115  ( .A(\normal/sll_15/n120 ), .B(
        \normal/sll_15/n112 ), .S0(n513), .Y(\normal/sll_15/n73 ) );
  MXI2X1 \normal/sll_15/U64  ( .A(\normal/sll_15/n77 ), .B(\normal/sll_15/n73 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n30 ) );
  MXI2X1 \normal/sll_15/U17  ( .A(\normal/sll_15/n31 ), .B(\normal/sll_15/n30 ), .S0(n503), .Y(\normal/N78 ) );
  MXI2X1 \normal/srl_15/U16  ( .A(\normal/srl_15/n32 ), .B(\normal/srl_15/n33 ), .S0(n503), .Y(\normal/N33 ) );
  MXI2X1 \normal/sll_15/U16  ( .A(\normal/sll_15/n32 ), .B(\normal/sll_15/n31 ), .S0(n503), .Y(\normal/N79 ) );
  MXI2X1 \normal/srl_15/U265  ( .A(\normal/srl_15/A[29] ), .B(add_out[45]), 
        .S0(n703), .Y(\normal/srl_15/n228 ) );
  MXI2X1 \normal/srl_15/U115  ( .A(\normal/srl_15/n128 ), .B(
        \normal/srl_15/n136 ), .S0(n513), .Y(\normal/srl_15/n78 ) );
  MXI2X1 \normal/srl_15/U65  ( .A(\normal/srl_15/n78 ), .B(\normal/srl_15/n82 ), .S0(n512), .Y(\normal/srl_15/n30 ) );
  MXI2X1 \normal/srl_15/U18  ( .A(\normal/srl_15/n30 ), .B(\normal/srl_15/n31 ), .S0(n503), .Y(\normal/N31 ) );
  MXI2X1 \normal/sll_15/U218  ( .A(\normal/sll_15/n205 ), .B(
        \normal/sll_15/n203 ), .S0(n514), .Y(\normal/sll_15/n158 ) );
  MXI2X1 \normal/sll_15/U116  ( .A(\normal/sll_15/n119 ), .B(
        \normal/sll_15/n111 ), .S0(n513), .Y(\normal/sll_15/n72 ) );
  MXI2X1 \normal/sll_15/U65  ( .A(\normal/sll_15/n76 ), .B(\normal/sll_15/n72 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n29 ) );
  MXI2X1 \normal/sll_15/U18  ( .A(\normal/sll_15/n30 ), .B(\normal/sll_15/n29 ), .S0(n503), .Y(\normal/N77 ) );
  MXI2X1 \normal/srl_15/U266  ( .A(add_out[28]), .B(\normal/srl_15/A[44] ), 
        .S0(n703), .Y(\normal/srl_15/n227 ) );
  MXI2X1 \normal/srl_15/U116  ( .A(\normal/srl_15/n127 ), .B(
        \normal/srl_15/n135 ), .S0(n513), .Y(\normal/srl_15/n77 ) );
  MXI2X1 \normal/srl_15/U66  ( .A(\normal/srl_15/n77 ), .B(\normal/srl_15/n81 ), .S0(n512), .Y(\normal/srl_15/n29 ) );
  MXI2X1 \normal/srl_15/U19  ( .A(\normal/srl_15/n29 ), .B(\normal/srl_15/n30 ), .S0(n503), .Y(\normal/N30 ) );
  MXI2X1 \normal/sll_15/U219  ( .A(\normal/sll_15/n204 ), .B(
        \normal/sll_15/n202 ), .S0(n514), .Y(\normal/sll_15/n157 ) );
  MXI2X1 \normal/sll_15/U117  ( .A(\normal/sll_15/n118 ), .B(
        \normal/sll_15/n110 ), .S0(n513), .Y(\normal/sll_15/n71 ) );
  MXI2X1 \normal/sll_15/U66  ( .A(\normal/sll_15/n75 ), .B(\normal/sll_15/n71 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n28 ) );
  MXI2X1 \normal/sll_15/U19  ( .A(\normal/sll_15/n29 ), .B(\normal/sll_15/n28 ), .S0(n503), .Y(\normal/N76 ) );
  MXI2X1 \normal/srl_15/U271  ( .A(add_out[23]), .B(add_out[39]), .S0(n714), 
        .Y(\normal/srl_15/n222 ) );
  MXI2X1 \normal/srl_15/U269  ( .A(\normal/srl_15/A[25] ), .B(
        \normal/srl_15/A[41] ), .S0(n714), .Y(\normal/srl_15/n224 ) );
  MXI2X1 \normal/srl_15/U121  ( .A(\normal/srl_15/n122 ), .B(
        \normal/srl_15/n130 ), .S0(n513), .Y(\normal/srl_15/n72 ) );
  MXI2X1 \normal/srl_15/U267  ( .A(\normal/srl_15/A[27] ), .B(add_out[43]), 
        .S0(n703), .Y(\normal/srl_15/n226 ) );
  MXI2X1 \normal/srl_15/U117  ( .A(\normal/srl_15/n126 ), .B(
        \normal/srl_15/n134 ), .S0(n513), .Y(\normal/srl_15/n76 ) );
  MXI2X1 \normal/srl_15/U270  ( .A(add_out[24]), .B(\normal/srl_15/A[40] ), 
        .S0(n714), .Y(\normal/srl_15/n223 ) );
  MXI2X1 \normal/srl_15/U268  ( .A(add_out[26]), .B(add_out[42]), .S0(n703), 
        .Y(\normal/srl_15/n225 ) );
  MXI2X1 \normal/srl_15/U220  ( .A(\normal/srl_15/n223 ), .B(
        \normal/srl_15/n225 ), .S0(n715), .Y(\normal/srl_15/n173 ) );
  MXI2X1 \normal/srl_15/U120  ( .A(\normal/srl_15/n123 ), .B(
        \normal/srl_15/n131 ), .S0(n513), .Y(\normal/srl_15/n73 ) );
  MXI2X1 \normal/srl_15/U70  ( .A(\normal/srl_15/n73 ), .B(\normal/srl_15/n77 ), .S0(n512), .Y(\normal/srl_15/n25 ) );
  MXI2X1 \normal/sll_15/U223  ( .A(\normal/sll_15/n200 ), .B(
        \normal/sll_15/n198 ), .S0(n514), .Y(\normal/sll_15/n153 ) );
  MXI2X1 \normal/sll_15/U121  ( .A(\normal/sll_15/n114 ), .B(
        \normal/sll_15/n106 ), .S0(n513), .Y(\normal/sll_15/n67 ) );
  MXI2X1 \normal/sll_15/U70  ( .A(\normal/sll_15/n71 ), .B(\normal/sll_15/n67 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n24 ) );
  MXI2X1 \normal/sll_15/U220  ( .A(\normal/sll_15/n203 ), .B(
        \normal/sll_15/n201 ), .S0(n514), .Y(\normal/sll_15/n156 ) );
  MXI2X1 \normal/sll_15/U118  ( .A(\normal/sll_15/n117 ), .B(
        \normal/sll_15/n109 ), .S0(n513), .Y(\normal/sll_15/n70 ) );
  MXI2X1 \normal/sll_15/U224  ( .A(\normal/sll_15/n199 ), .B(
        \normal/sll_15/n197 ), .S0(n514), .Y(\normal/sll_15/n152 ) );
  MXI2X1 \normal/sll_15/U122  ( .A(\normal/sll_15/n113 ), .B(
        \normal/sll_15/n105 ), .S0(n513), .Y(\normal/sll_15/n66 ) );
  MXI2X1 \normal/srl_15/U219  ( .A(\normal/srl_15/n224 ), .B(
        \normal/srl_15/n226 ), .S0(n715), .Y(\normal/srl_15/n174 ) );
  MXI2X1 \normal/srl_15/U119  ( .A(\normal/srl_15/n124 ), .B(
        \normal/srl_15/n132 ), .S0(n513), .Y(\normal/srl_15/n74 ) );
  MXI2X1 \normal/srl_15/U69  ( .A(\normal/srl_15/n74 ), .B(\normal/srl_15/n78 ), .S0(n704), .Y(\normal/srl_15/n26 ) );
  MXI2X1 \normal/srl_15/U23  ( .A(\normal/srl_15/n25 ), .B(\normal/srl_15/n26 ), .S0(n503), .Y(\normal/N26 ) );
  MXI2X1 \normal/sll_15/U222  ( .A(\normal/sll_15/n201 ), .B(
        \normal/sll_15/n199 ), .S0(n514), .Y(\normal/sll_15/n154 ) );
  MXI2X1 \normal/sll_15/U120  ( .A(\normal/sll_15/n115 ), .B(
        \normal/sll_15/n107 ), .S0(n513), .Y(\normal/sll_15/n68 ) );
  MXI2X1 \normal/sll_15/U69  ( .A(\normal/sll_15/n72 ), .B(\normal/sll_15/n68 ), .S0(n704), .Y(\normal/sll_15/n25 ) );
  MXI2X1 \normal/sll_15/U23  ( .A(\normal/sll_15/n25 ), .B(\normal/sll_15/n24 ), .S0(n503), .Y(\normal/N72 ) );
  MXI2X1 \normal/srl_15/U218  ( .A(\normal/srl_15/n225 ), .B(
        \normal/srl_15/n227 ), .S0(n715), .Y(\normal/srl_15/n175 ) );
  MXI2X1 \normal/srl_15/U118  ( .A(\normal/srl_15/n125 ), .B(
        \normal/srl_15/n133 ), .S0(n513), .Y(\normal/srl_15/n75 ) );
  MXI2X1 \normal/srl_15/U68  ( .A(\normal/srl_15/n75 ), .B(\normal/srl_15/n79 ), .S0(n512), .Y(\normal/srl_15/n27 ) );
  MXI2X1 \normal/srl_15/U22  ( .A(\normal/srl_15/n26 ), .B(\normal/srl_15/n27 ), .S0(n503), .Y(\normal/N27 ) );
  MXI2X1 \normal/sll_15/U221  ( .A(\normal/sll_15/n202 ), .B(
        \normal/sll_15/n200 ), .S0(n514), .Y(\normal/sll_15/n155 ) );
  MXI2X1 \normal/sll_15/U119  ( .A(\normal/sll_15/n116 ), .B(
        \normal/sll_15/n108 ), .S0(n513), .Y(\normal/sll_15/n69 ) );
  MXI2X1 \normal/sll_15/U68  ( .A(\normal/sll_15/n73 ), .B(\normal/sll_15/n69 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n26 ) );
  MXI2X1 \normal/sll_15/U22  ( .A(\normal/sll_15/n26 ), .B(\normal/sll_15/n25 ), .S0(n503), .Y(\normal/N73 ) );
  MXI2X1 \normal/srl_15/U67  ( .A(\normal/srl_15/n76 ), .B(\normal/srl_15/n80 ), .S0(n512), .Y(\normal/srl_15/n28 ) );
  MXI2X1 \normal/sll_15/U67  ( .A(\normal/sll_15/n74 ), .B(\normal/sll_15/n70 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n27 ) );
  MXI2X1 \normal/srl_15/U21  ( .A(\normal/srl_15/n27 ), .B(\normal/srl_15/n28 ), .S0(n503), .Y(\normal/N28 ) );
  MXI2X1 \normal/sll_15/U21  ( .A(\normal/sll_15/n27 ), .B(\normal/sll_15/n26 ), .S0(n503), .Y(\normal/N74 ) );
  MXI2X1 \normal/srl_15/U49  ( .A(\normal/srl_15/n94 ), .B(\normal/srl_15/n98 ), .S0(n704), .Y(\normal/srl_15/n46 ) );
  MXI2X1 \normal/sll_15/U238  ( .A(add_out[43]), .B(\normal/srl_15/A[27] ), 
        .S0(n703), .Y(\normal/sll_15/n232 ) );
  MXI2X1 \normal/sll_15/U142  ( .A(\normal/sll_15/n187 ), .B(
        \normal/sll_15/n155 ), .S0(n504), .Y(\normal/sll_15/n140 ) );
  MXI2X1 \normal/sll_15/U95  ( .A(\normal/sll_15/n140 ), .B(
        \normal/sll_15/n132 ), .S0(n513), .Y(\normal/sll_15/n93 ) );
  MXI2X1 \normal/sll_15/U240  ( .A(\normal/srl_15/A[41] ), .B(
        \normal/srl_15/A[25] ), .S0(n703), .Y(\normal/sll_15/n230 ) );
  MXI2X1 \normal/sll_15/U193  ( .A(\normal/sll_15/n230 ), .B(
        \normal/sll_15/n228 ), .S0(n514), .Y(\normal/sll_15/n183 ) );
  MXI2X1 \normal/sll_15/U225  ( .A(\normal/sll_15/n198 ), .B(
        \normal/sll_15/n196 ), .S0(n514), .Y(\normal/sll_15/n151 ) );
  MXI2X1 \normal/sll_15/U146  ( .A(\normal/sll_15/n183 ), .B(
        \normal/sll_15/n151 ), .S0(n504), .Y(\normal/sll_15/n136 ) );
  MXI2X1 \normal/sll_15/U99  ( .A(\normal/sll_15/n136 ), .B(
        \normal/sll_15/n128 ), .S0(n513), .Y(\normal/sll_15/n89 ) );
  MXI2X1 \normal/sll_15/U237  ( .A(\normal/srl_15/A[44] ), .B(add_out[28]), 
        .S0(n714), .Y(\normal/sll_15/n233 ) );
  MXI2X1 \normal/sll_15/U239  ( .A(add_out[42]), .B(add_out[26]), .S0(n703), 
        .Y(\normal/sll_15/n231 ) );
  MXI2X1 \normal/sll_15/U143  ( .A(\normal/sll_15/n186 ), .B(
        \normal/sll_15/n154 ), .S0(n504), .Y(\normal/sll_15/n139 ) );
  MXI2X1 \normal/sll_15/U96  ( .A(\normal/sll_15/n139 ), .B(
        \normal/sll_15/n131 ), .S0(n513), .Y(\normal/sll_15/n92 ) );
  MXI2X1 \normal/sll_15/U241  ( .A(\normal/srl_15/A[40] ), .B(add_out[24]), 
        .S0(n703), .Y(\normal/sll_15/n229 ) );
  MXI2X1 \normal/sll_15/U194  ( .A(\normal/sll_15/n229 ), .B(
        \normal/sll_15/n227 ), .S0(n514), .Y(\normal/sll_15/n182 ) );
  MXI2X1 \normal/sll_15/U226  ( .A(\normal/sll_15/n197 ), .B(
        \normal/sll_15/n195 ), .S0(n514), .Y(\normal/sll_15/n150 ) );
  MXI2X1 \normal/sll_15/U147  ( .A(\normal/sll_15/n182 ), .B(
        \normal/sll_15/n150 ), .S0(n504), .Y(\normal/sll_15/n135 ) );
  MXI2X1 \normal/sll_15/U100  ( .A(\normal/sll_15/n135 ), .B(
        \normal/sll_15/n127 ), .S0(n513), .Y(\normal/sll_15/n88 ) );
  MXI2X1 \normal/srl_15/U50  ( .A(\normal/srl_15/n93 ), .B(\normal/srl_15/n97 ), .S0(n704), .Y(\normal/srl_15/n45 ) );
  MXI2X1 \normal/sll_15/U144  ( .A(\normal/sll_15/n185 ), .B(
        \normal/sll_15/n153 ), .S0(n504), .Y(\normal/sll_15/n138 ) );
  MXI2X1 \normal/sll_15/U97  ( .A(\normal/sll_15/n138 ), .B(
        \normal/sll_15/n130 ), .S0(n513), .Y(\normal/sll_15/n91 ) );
  MXI2X1 \normal/srl_15/U1  ( .A(\normal/srl_15/n47 ), .B(\normal/srl_15/n48 ), 
        .S0(n503), .Y(\normal/N48 ) );
  MXI2X1 \normal/sll_15/U141  ( .A(\normal/sll_15/n188 ), .B(
        \normal/sll_15/n156 ), .S0(n504), .Y(\normal/sll_15/n141 ) );
  MXI2X1 \normal/sll_15/U94  ( .A(\normal/sll_15/n141 ), .B(
        \normal/sll_15/n133 ), .S0(n513), .Y(\normal/sll_15/n94 ) );
  MXI2X1 \normal/sll_15/U192  ( .A(\normal/sll_15/n231 ), .B(
        \normal/sll_15/n229 ), .S0(n514), .Y(\normal/sll_15/n184 ) );
  MXI2X1 \normal/sll_15/U145  ( .A(\normal/sll_15/n184 ), .B(
        \normal/sll_15/n152 ), .S0(n504), .Y(\normal/sll_15/n137 ) );
  MXI2X1 \normal/sll_15/U98  ( .A(\normal/sll_15/n137 ), .B(
        \normal/sll_15/n129 ), .S0(n513), .Y(\normal/sll_15/n90 ) );
  MXI2X1 \normal/sll_15/U47  ( .A(\normal/sll_15/n94 ), .B(\normal/sll_15/n90 ), .S0(n704), .Y(\normal/sll_15/n47 ) );
  MXI2X1 \normal/srl_15/U53  ( .A(\normal/srl_15/n90 ), .B(\normal/srl_15/n94 ), .S0(n704), .Y(\normal/srl_15/n42 ) );
  MXI2X1 \normal/srl_15/U52  ( .A(\normal/srl_15/n91 ), .B(\normal/srl_15/n95 ), .S0(n704), .Y(\normal/srl_15/n43 ) );
  MXI2X1 \normal/srl_15/U6  ( .A(\normal/srl_15/n42 ), .B(\normal/srl_15/n43 ), 
        .S0(n503), .Y(\normal/N43 ) );
  MXI2X1 \normal/sll_15/U6  ( .A(\normal/sll_15/n42 ), .B(\normal/sll_15/n41 ), 
        .S0(n503), .Y(\normal/N89 ) );
  MXI2X1 \normal/srl_15/U7  ( .A(\normal/srl_15/n41 ), .B(\normal/srl_15/n42 ), 
        .S0(n503), .Y(\normal/N42 ) );
  MXI2X1 \normal/srl_15/U51  ( .A(\normal/srl_15/n92 ), .B(\normal/srl_15/n96 ), .S0(n704), .Y(\normal/srl_15/n44 ) );
  MXI2X1 \normal/srl_15/U5  ( .A(\normal/srl_15/n43 ), .B(\normal/srl_15/n44 ), 
        .S0(n503), .Y(\normal/N44 ) );
  MXI2X1 \normal/sll_15/U5  ( .A(\normal/sll_15/n43 ), .B(\normal/sll_15/n42 ), 
        .S0(n503), .Y(\normal/N90 ) );
  MXI2X1 \normal/srl_15/U4  ( .A(\normal/srl_15/n44 ), .B(\normal/srl_15/n45 ), 
        .S0(n503), .Y(\normal/N45 ) );
  MXI2X1 \normal/sll_15/U4  ( .A(\normal/sll_15/n44 ), .B(\normal/sll_15/n43 ), 
        .S0(n503), .Y(\normal/N91 ) );
  MXI2X1 \normal/srl_15/U291  ( .A(add_out[3]), .B(add_out[19]), .S0(n703), 
        .Y(\normal/srl_15/n202 ) );
  MXI2X1 \normal/srl_15/U285  ( .A(\normal/srl_15/A[9] ), .B(
        \normal/srl_15/A[25] ), .S0(n703), .Y(\normal/srl_15/n208 ) );
  MXI2X1 \normal/srl_15/U283  ( .A(\normal/srl_15/A[11] ), .B(
        \normal/srl_15/A[27] ), .S0(n703), .Y(\normal/srl_15/n210 ) );
  MXI2X1 \normal/srl_15/U185  ( .A(\normal/srl_15/n158 ), .B(
        \normal/srl_15/n190 ), .S0(n504), .Y(\normal/srl_15/n108 ) );
  MXI2X1 \normal/srl_15/U143  ( .A(\normal/srl_15/n100 ), .B(
        \normal/srl_15/n108 ), .S0(n513), .Y(\normal/srl_15/n50 ) );
  MXI2X1 \normal/srl_15/U289  ( .A(add_out[5]), .B(\normal/srl_15/A[21] ), 
        .S0(n703), .Y(\normal/srl_15/n204 ) );
  MXI2X1 \normal/srl_15/U287  ( .A(add_out[7]), .B(add_out[23]), .S0(n703), 
        .Y(\normal/srl_15/n206 ) );
  MXI2X1 \normal/srl_15/U189  ( .A(\normal/srl_15/n154 ), .B(
        \normal/srl_15/n186 ), .S0(n504), .Y(\normal/srl_15/n104 ) );
  MXI2X1 \normal/srl_15/U281  ( .A(add_out[13]), .B(\normal/srl_15/A[29] ), 
        .S0(n714), .Y(\normal/srl_15/n212 ) );
  MXI2X1 \normal/srl_15/U279  ( .A(add_out[15]), .B(add_out[31]), .S0(n714), 
        .Y(\normal/srl_15/n214 ) );
  MXI2X1 \normal/srl_15/U231  ( .A(\normal/srl_15/n212 ), .B(
        \normal/srl_15/n214 ), .S0(n715), .Y(\normal/srl_15/n162 ) );
  MXI2X1 \normal/srl_15/U181  ( .A(\normal/srl_15/n162 ), .B(
        \normal/srl_15/n194 ), .S0(n504), .Y(\normal/srl_15/n112 ) );
  MXI2X1 \normal/srl_15/U139  ( .A(\normal/srl_15/n104 ), .B(
        \normal/srl_15/n112 ), .S0(n513), .Y(\normal/srl_15/n54 ) );
  MXI2X1 \normal/srl_15/U93  ( .A(\normal/srl_15/n50 ), .B(\normal/srl_15/n54 ), .S0(n512), .Y(\normal/srl_15/n2 ) );
  MXI2X1 \normal/srl_15/U292  ( .A(add_out[2]), .B(add_out[18]), .S0(n703), 
        .Y(\normal/srl_15/n201 ) );
  MXI2X1 \normal/srl_15/U290  ( .A(\normal/srl_15/A[4] ), .B(add_out[20]), 
        .S0(n703), .Y(\normal/srl_15/n203 ) );
  MXI2X1 \normal/srl_15/U284  ( .A(\normal/srl_15/A[10] ), .B(add_out[26]), 
        .S0(n703), .Y(\normal/srl_15/n209 ) );
  MXI2X1 \normal/srl_15/U282  ( .A(\normal/srl_15/A[12] ), .B(add_out[28]), 
        .S0(n703), .Y(\normal/srl_15/n211 ) );
  MXI2X1 \normal/srl_15/U184  ( .A(\normal/srl_15/n159 ), .B(
        \normal/srl_15/n191 ), .S0(n504), .Y(\normal/srl_15/n109 ) );
  MXI2X1 \normal/srl_15/U142  ( .A(\normal/srl_15/n101 ), .B(
        \normal/srl_15/n109 ), .S0(n513), .Y(\normal/srl_15/n51 ) );
  MXI2X1 \normal/srl_15/U288  ( .A(\normal/srl_15/A[6] ), .B(
        \normal/srl_15/A[22] ), .S0(n703), .Y(\normal/srl_15/n205 ) );
  MXI2X1 \normal/srl_15/U286  ( .A(\normal/srl_15/A[8] ), .B(add_out[24]), 
        .S0(n703), .Y(\normal/srl_15/n207 ) );
  MXI2X1 \normal/srl_15/U188  ( .A(\normal/srl_15/n155 ), .B(
        \normal/srl_15/n187 ), .S0(n504), .Y(\normal/srl_15/n105 ) );
  MXI2X1 \normal/srl_15/U280  ( .A(add_out[14]), .B(add_out[30]), .S0(n714), 
        .Y(\normal/srl_15/n213 ) );
  MXI2X1 \normal/srl_15/U278  ( .A(add_out[16]), .B(\normal/srl_15/A[32] ), 
        .S0(n714), .Y(\normal/srl_15/n215 ) );
  MXI2X1 \normal/srl_15/U230  ( .A(\normal/srl_15/n213 ), .B(
        \normal/srl_15/n215 ), .S0(n715), .Y(\normal/srl_15/n163 ) );
  MXI2X1 \normal/srl_15/U180  ( .A(\normal/srl_15/n163 ), .B(
        \normal/srl_15/n195 ), .S0(n504), .Y(\normal/srl_15/n113 ) );
  MXI2X1 \normal/srl_15/U138  ( .A(\normal/srl_15/n105 ), .B(
        \normal/srl_15/n113 ), .S0(n513), .Y(\normal/srl_15/n55 ) );
  MXI2X1 \normal/srl_15/U92  ( .A(\normal/srl_15/n51 ), .B(\normal/srl_15/n55 ), .S0(n512), .Y(\normal/srl_15/n3 ) );
  MXI2X1 \normal/srl_15/U45  ( .A(\normal/srl_15/n2 ), .B(\normal/srl_15/n3 ), 
        .S0(n503), .Y(\normal/N4 ) );
  MXI2X1 \normal/srl_15/U183  ( .A(\normal/srl_15/n160 ), .B(
        \normal/srl_15/n192 ), .S0(n504), .Y(\normal/srl_15/n110 ) );
  MXI2X1 \normal/srl_15/U141  ( .A(\normal/srl_15/n102 ), .B(
        \normal/srl_15/n110 ), .S0(n513), .Y(\normal/srl_15/n52 ) );
  MXI2X1 \normal/srl_15/U187  ( .A(\normal/srl_15/n156 ), .B(
        \normal/srl_15/n188 ), .S0(n504), .Y(\normal/srl_15/n106 ) );
  MXI2X1 \normal/srl_15/U277  ( .A(add_out[17]), .B(add_out[33]), .S0(n714), 
        .Y(\normal/srl_15/n216 ) );
  MXI2X1 \normal/srl_15/U229  ( .A(\normal/srl_15/n214 ), .B(
        \normal/srl_15/n216 ), .S0(n715), .Y(\normal/srl_15/n164 ) );
  MXI2X1 \normal/srl_15/U179  ( .A(\normal/srl_15/n164 ), .B(
        \normal/srl_15/n196 ), .S0(n504), .Y(\normal/srl_15/n114 ) );
  MXI2X1 \normal/srl_15/U137  ( .A(\normal/srl_15/n106 ), .B(
        \normal/srl_15/n114 ), .S0(n513), .Y(\normal/srl_15/n56 ) );
  MXI2X1 \normal/srl_15/U91  ( .A(\normal/srl_15/n52 ), .B(\normal/srl_15/n56 ), .S0(n512), .Y(\normal/srl_15/n4 ) );
  MXI2X1 \normal/srl_15/U44  ( .A(\normal/srl_15/n3 ), .B(\normal/srl_15/n4 ), 
        .S0(n503), .Y(\normal/N5 ) );
  MXI2X1 \normal/srl_15/U190  ( .A(\normal/srl_15/n153 ), .B(
        \normal/srl_15/n185 ), .S0(n504), .Y(\normal/srl_15/n103 ) );
  MXI2X1 \normal/srl_15/U182  ( .A(\normal/srl_15/n161 ), .B(
        \normal/srl_15/n193 ), .S0(n504), .Y(\normal/srl_15/n111 ) );
  MXI2X1 \normal/srl_15/U140  ( .A(\normal/srl_15/n103 ), .B(
        \normal/srl_15/n111 ), .S0(n513), .Y(\normal/srl_15/n53 ) );
  MXI2X1 \normal/srl_15/U186  ( .A(\normal/srl_15/n157 ), .B(
        \normal/srl_15/n189 ), .S0(n504), .Y(\normal/srl_15/n107 ) );
  MXI2X1 \normal/srl_15/U276  ( .A(add_out[18]), .B(add_out[34]), .S0(n714), 
        .Y(\normal/srl_15/n217 ) );
  MXI2X1 \normal/srl_15/U228  ( .A(\normal/srl_15/n215 ), .B(
        \normal/srl_15/n217 ), .S0(n715), .Y(\normal/srl_15/n165 ) );
  MXI2X1 \normal/srl_15/U178  ( .A(\normal/srl_15/n165 ), .B(
        \normal/srl_15/n197 ), .S0(n504), .Y(\normal/srl_15/n115 ) );
  MXI2X1 \normal/srl_15/U136  ( .A(\normal/srl_15/n107 ), .B(
        \normal/srl_15/n115 ), .S0(n513), .Y(\normal/srl_15/n57 ) );
  MXI2X1 \normal/srl_15/U90  ( .A(\normal/srl_15/n53 ), .B(\normal/srl_15/n57 ), .S0(n512), .Y(\normal/srl_15/n5 ) );
  MXI2X1 \normal/srl_15/U43  ( .A(\normal/srl_15/n4 ), .B(\normal/srl_15/n5 ), 
        .S0(n503), .Y(\normal/N6 ) );
  MXI2X1 \normal/srl_15/U275  ( .A(add_out[19]), .B(add_out[35]), .S0(n714), 
        .Y(\normal/srl_15/n218 ) );
  MXI2X1 \normal/srl_15/U227  ( .A(\normal/srl_15/n216 ), .B(
        \normal/srl_15/n218 ), .S0(n715), .Y(\normal/srl_15/n166 ) );
  MXI2X1 \normal/srl_15/U177  ( .A(\normal/srl_15/n166 ), .B(
        \normal/srl_15/n198 ), .S0(n504), .Y(\normal/srl_15/n116 ) );
  MXI2X1 \normal/srl_15/U135  ( .A(\normal/srl_15/n108 ), .B(
        \normal/srl_15/n116 ), .S0(n513), .Y(\normal/srl_15/n58 ) );
  MXI2X1 \normal/srl_15/U89  ( .A(\normal/srl_15/n54 ), .B(\normal/srl_15/n58 ), .S0(n512), .Y(\normal/srl_15/n6 ) );
  MXI2X1 \normal/srl_15/U42  ( .A(\normal/srl_15/n5 ), .B(\normal/srl_15/n6 ), 
        .S0(n503), .Y(\normal/N7 ) );
  MXI2X1 \normal/srl_15/U274  ( .A(add_out[20]), .B(\normal/srl_15/A[36] ), 
        .S0(n714), .Y(\normal/srl_15/n219 ) );
  MXI2X1 \normal/srl_15/U134  ( .A(\normal/srl_15/n109 ), .B(
        \normal/srl_15/n117 ), .S0(n513), .Y(\normal/srl_15/n59 ) );
  MXI2X1 \normal/srl_15/U88  ( .A(\normal/srl_15/n55 ), .B(\normal/srl_15/n59 ), .S0(n512), .Y(\normal/srl_15/n7 ) );
  MXI2X1 \normal/srl_15/U41  ( .A(\normal/srl_15/n6 ), .B(\normal/srl_15/n7 ), 
        .S0(n503), .Y(\normal/N8 ) );
  MXI2X1 \normal/srl_15/U273  ( .A(\normal/srl_15/A[21] ), .B(add_out[37]), 
        .S0(n714), .Y(\normal/srl_15/n220 ) );
  MXI2X1 \normal/srl_15/U133  ( .A(\normal/srl_15/n110 ), .B(
        \normal/srl_15/n118 ), .S0(n513), .Y(\normal/srl_15/n60 ) );
  MXI2X1 \normal/srl_15/U87  ( .A(\normal/srl_15/n56 ), .B(\normal/srl_15/n60 ), .S0(n512), .Y(\normal/srl_15/n8 ) );
  MXI2X1 \normal/srl_15/U40  ( .A(\normal/srl_15/n7 ), .B(\normal/srl_15/n8 ), 
        .S0(n503), .Y(\normal/N9 ) );
  MXI2X1 \normal/srl_15/U272  ( .A(\normal/srl_15/A[22] ), .B(add_out[38]), 
        .S0(n714), .Y(\normal/srl_15/n221 ) );
  MXI2X1 \normal/srl_15/U224  ( .A(\normal/srl_15/n219 ), .B(
        \normal/srl_15/n221 ), .S0(n715), .Y(\normal/srl_15/n169 ) );
  MXI2X1 \normal/srl_15/U132  ( .A(\normal/srl_15/n111 ), .B(
        \normal/srl_15/n119 ), .S0(n513), .Y(\normal/srl_15/n61 ) );
  MXI2X1 \normal/srl_15/U86  ( .A(\normal/srl_15/n57 ), .B(\normal/srl_15/n61 ), .S0(n512), .Y(\normal/srl_15/n9 ) );
  MXI2X1 \normal/srl_15/U39  ( .A(\normal/srl_15/n8 ), .B(\normal/srl_15/n9 ), 
        .S0(n503), .Y(\normal/N10 ) );
  MXI2X1 \normal/srl_15/U131  ( .A(\normal/srl_15/n112 ), .B(
        \normal/srl_15/n120 ), .S0(n513), .Y(\normal/srl_15/n62 ) );
  MXI2X1 \normal/srl_15/U85  ( .A(\normal/srl_15/n58 ), .B(\normal/srl_15/n62 ), .S0(n512), .Y(\normal/srl_15/n10 ) );
  MXI2X1 \normal/srl_15/U38  ( .A(\normal/srl_15/n9 ), .B(\normal/srl_15/n10 ), 
        .S0(n503), .Y(\normal/N11 ) );
  MXI2X1 \normal/srl_15/U127  ( .A(\normal/srl_15/n116 ), .B(
        \normal/srl_15/n124 ), .S0(n513), .Y(\normal/srl_15/n66 ) );
  MXI2X1 \normal/srl_15/U123  ( .A(\normal/srl_15/n120 ), .B(
        \normal/srl_15/n128 ), .S0(n513), .Y(\normal/srl_15/n70 ) );
  MXI2X1 \normal/srl_15/U77  ( .A(\normal/srl_15/n66 ), .B(\normal/srl_15/n70 ), .S0(n704), .Y(\normal/srl_15/n18 ) );
  MXI2X1 \normal/srl_15/U126  ( .A(\normal/srl_15/n117 ), .B(
        \normal/srl_15/n125 ), .S0(n513), .Y(\normal/srl_15/n67 ) );
  MXI2X1 \normal/srl_15/U122  ( .A(\normal/srl_15/n121 ), .B(
        \normal/srl_15/n129 ), .S0(n513), .Y(\normal/srl_15/n71 ) );
  MXI2X1 \normal/srl_15/U76  ( .A(\normal/srl_15/n67 ), .B(\normal/srl_15/n71 ), .S0(n704), .Y(\normal/srl_15/n19 ) );
  MXI2X1 \normal/srl_15/U125  ( .A(\normal/srl_15/n118 ), .B(
        \normal/srl_15/n126 ), .S0(n513), .Y(\normal/srl_15/n68 ) );
  MXI2X1 \normal/srl_15/U75  ( .A(\normal/srl_15/n68 ), .B(\normal/srl_15/n72 ), .S0(n704), .Y(\normal/srl_15/n20 ) );
  MXI2X1 \normal/srl_15/U73  ( .A(\normal/srl_15/n70 ), .B(\normal/srl_15/n74 ), .S0(n704), .Y(\normal/srl_15/n22 ) );
  MXI2X1 \normal/srl_15/U26  ( .A(\normal/srl_15/n22 ), .B(\normal/srl_15/n23 ), .S0(n503), .Y(\normal/N23 ) );
  MXI2X1 \normal/srl_15/U144  ( .A(\normal/srl_15/n99 ), .B(
        \normal/srl_15/n107 ), .S0(n513), .Y(\normal/srl_15/n49 ) );
  MXI2X1 \normal/srl_15/U94  ( .A(\normal/srl_15/n49 ), .B(\normal/srl_15/n53 ), .S0(n512), .Y(\normal/srl_15/n1 ) );
  MXI2X1 \normal/srl_15/U46  ( .A(\normal/srl_15/n1 ), .B(\normal/srl_15/n2 ), 
        .S0(n503), .Y(\normal/N3 ) );
  MXI2X1 \normal/srl_15/U124  ( .A(\normal/srl_15/n119 ), .B(
        \normal/srl_15/n127 ), .S0(n513), .Y(\normal/srl_15/n69 ) );
  MXI2X1 \normal/srl_15/U74  ( .A(\normal/srl_15/n69 ), .B(\normal/srl_15/n73 ), .S0(n704), .Y(\normal/srl_15/n21 ) );
  MXI2X1 \normal/srl_15/U27  ( .A(\normal/srl_15/n20 ), .B(\normal/srl_15/n21 ), .S0(n503), .Y(\normal/N22 ) );
  MXI2X1 \normal/srl_15/U130  ( .A(\normal/srl_15/n113 ), .B(
        \normal/srl_15/n121 ), .S0(n513), .Y(\normal/srl_15/n63 ) );
  MXI2X1 \normal/srl_15/U84  ( .A(\normal/srl_15/n59 ), .B(\normal/srl_15/n63 ), .S0(n512), .Y(\normal/srl_15/n11 ) );
  MXI2X1 \normal/srl_15/U129  ( .A(\normal/srl_15/n114 ), .B(
        \normal/srl_15/n122 ), .S0(n513), .Y(\normal/srl_15/n64 ) );
  MXI2X1 \normal/srl_15/U83  ( .A(\normal/srl_15/n60 ), .B(\normal/srl_15/n64 ), .S0(n512), .Y(\normal/srl_15/n12 ) );
  MXI2X1 \normal/srl_15/U128  ( .A(\normal/srl_15/n115 ), .B(
        \normal/srl_15/n123 ), .S0(n513), .Y(\normal/srl_15/n65 ) );
  MXI2X1 \normal/srl_15/U82  ( .A(\normal/srl_15/n61 ), .B(\normal/srl_15/n65 ), .S0(n512), .Y(\normal/srl_15/n13 ) );
  MXI2X1 \normal/srl_15/U35  ( .A(\normal/srl_15/n12 ), .B(\normal/srl_15/n13 ), .S0(n503), .Y(\normal/N14 ) );
  MXI2X1 \normal/srl_15/U81  ( .A(\normal/srl_15/n62 ), .B(\normal/srl_15/n66 ), .S0(n704), .Y(\normal/srl_15/n14 ) );
  MXI2X1 \normal/srl_15/U34  ( .A(\normal/srl_15/n13 ), .B(\normal/srl_15/n14 ), .S0(n503), .Y(\normal/N15 ) );
  MXI2X1 \normal/srl_15/U80  ( .A(\normal/srl_15/n63 ), .B(\normal/srl_15/n67 ), .S0(n704), .Y(\normal/srl_15/n15 ) );
  MXI2X1 \normal/srl_15/U79  ( .A(\normal/srl_15/n64 ), .B(\normal/srl_15/n68 ), .S0(n704), .Y(\normal/srl_15/n16 ) );
  MXI2X1 \normal/srl_15/U78  ( .A(\normal/srl_15/n65 ), .B(\normal/srl_15/n69 ), .S0(n704), .Y(\normal/srl_15/n17 ) );
  MXI2X1 \normal/sll_15/U131  ( .A(\normal/sll_15/n104 ), .B(
        \normal/sll_15/n96 ), .S0(n513), .Y(\normal/sll_15/n57 ) );
  MXI2X1 \normal/sll_15/U84  ( .A(\normal/sll_15/n57 ), .B(\normal/sll_15/n53 ), .S0(n512), .Y(\normal/sll_15/n10 ) );
  MXI2X1 \normal/sll_15/U132  ( .A(\normal/sll_15/n103 ), .B(
        \normal/sll_15/n95 ), .S0(n513), .Y(\normal/sll_15/n56 ) );
  MXI2X1 \normal/sll_15/U85  ( .A(\normal/sll_15/n56 ), .B(\normal/sll_15/n52 ), .S0(n512), .Y(\normal/sll_15/n9 ) );
  MXI2X1 \normal/sll_15/U37  ( .A(\normal/sll_15/n10 ), .B(\normal/sll_15/n9 ), 
        .S0(n503), .Y(\normal/N58 ) );
  MXI2X1 \normal/sll_15/U130  ( .A(\normal/sll_15/n105 ), .B(
        \normal/sll_15/n97 ), .S0(n513), .Y(\normal/sll_15/n58 ) );
  MXI2X1 \normal/sll_15/U83  ( .A(\normal/sll_15/n58 ), .B(\normal/sll_15/n54 ), .S0(n512), .Y(\normal/sll_15/n11 ) );
  MXI2X1 \normal/sll_15/U36  ( .A(\normal/sll_15/n11 ), .B(\normal/sll_15/n10 ), .S0(n503), .Y(\normal/N59 ) );
  MXI2X1 \normal/sll_15/U129  ( .A(\normal/sll_15/n106 ), .B(
        \normal/sll_15/n98 ), .S0(n513), .Y(\normal/sll_15/n59 ) );
  MXI2X1 \normal/sll_15/U82  ( .A(\normal/sll_15/n59 ), .B(\normal/sll_15/n55 ), .S0(n512), .Y(\normal/sll_15/n12 ) );
  MXI2X1 \normal/sll_15/U35  ( .A(\normal/sll_15/n12 ), .B(\normal/sll_15/n11 ), .S0(n503), .Y(\normal/N60 ) );
  MXI2X1 \normal/sll_15/U128  ( .A(\normal/sll_15/n107 ), .B(
        \normal/sll_15/n99 ), .S0(n513), .Y(\normal/sll_15/n60 ) );
  MXI2X1 \normal/sll_15/U81  ( .A(\normal/sll_15/n60 ), .B(\normal/sll_15/n56 ), .S0(n512), .Y(\normal/sll_15/n13 ) );
  MXI2X1 \normal/sll_15/U34  ( .A(\normal/sll_15/n13 ), .B(\normal/sll_15/n12 ), .S0(n503), .Y(\normal/N61 ) );
  MXI2X1 \normal/sll_15/U127  ( .A(\normal/sll_15/n108 ), .B(
        \normal/sll_15/n100 ), .S0(n513), .Y(\normal/sll_15/n61 ) );
  MXI2X1 \normal/sll_15/U80  ( .A(\normal/sll_15/n61 ), .B(\normal/sll_15/n57 ), .S0(n512), .Y(\normal/sll_15/n14 ) );
  MXI2X1 \normal/sll_15/U33  ( .A(\normal/sll_15/n14 ), .B(\normal/sll_15/n13 ), .S0(n503), .Y(\normal/N62 ) );
  MXI2X1 \normal/sll_15/U126  ( .A(\normal/sll_15/n109 ), .B(
        \normal/sll_15/n101 ), .S0(n513), .Y(\normal/sll_15/n62 ) );
  MXI2X1 \normal/sll_15/U79  ( .A(\normal/sll_15/n62 ), .B(\normal/sll_15/n58 ), .S0(n512), .Y(\normal/sll_15/n15 ) );
  MXI2X1 \normal/sll_15/U32  ( .A(\normal/sll_15/n15 ), .B(\normal/sll_15/n14 ), .S0(n503), .Y(\normal/N63 ) );
  MXI2X1 \normal/sll_15/U125  ( .A(\normal/sll_15/n110 ), .B(
        \normal/sll_15/n102 ), .S0(n513), .Y(\normal/sll_15/n63 ) );
  MXI2X1 \normal/sll_15/U78  ( .A(\normal/sll_15/n63 ), .B(\normal/sll_15/n59 ), .S0(n512), .Y(\normal/sll_15/n16 ) );
  MXI2X1 \normal/sll_15/U31  ( .A(\normal/sll_15/n16 ), .B(\normal/sll_15/n15 ), .S0(n503), .Y(\normal/N64 ) );
  MXI2X1 \normal/sll_15/U124  ( .A(\normal/sll_15/n111 ), .B(
        \normal/sll_15/n103 ), .S0(n513), .Y(\normal/sll_15/n64 ) );
  MXI2X1 \normal/sll_15/U77  ( .A(\normal/sll_15/n64 ), .B(\normal/sll_15/n60 ), .S0(n512), .Y(\normal/sll_15/n17 ) );
  MXI2X1 \normal/sll_15/U30  ( .A(\normal/sll_15/n17 ), .B(\normal/sll_15/n16 ), .S0(n503), .Y(\normal/N65 ) );
  MXI2X1 \normal/sll_15/U89  ( .A(\normal/sll_15/n52 ), .B(\normal/sll_15/n48 ), .S0(n704), .Y(\normal/sll_15/n5 ) );
  MXI2X1 \normal/sll_15/U74  ( .A(\normal/sll_15/n67 ), .B(\normal/sll_15/n63 ), .S0(n512), .Y(\normal/sll_15/n20 ) );
  MXI2X1 \normal/sll_15/U75  ( .A(\normal/sll_15/n66 ), .B(\normal/sll_15/n62 ), .S0(n512), .Y(\normal/sll_15/n19 ) );
  MXI2X1 \normal/sll_15/U27  ( .A(\normal/sll_15/n20 ), .B(\normal/sll_15/n19 ), .S0(n503), .Y(\normal/N68 ) );
  MXI2X1 \normal/sll_15/U123  ( .A(\normal/sll_15/n112 ), .B(
        \normal/sll_15/n104 ), .S0(n513), .Y(\normal/sll_15/n65 ) );
  MXI2X1 \normal/sll_15/U73  ( .A(\normal/sll_15/n68 ), .B(\normal/sll_15/n64 ), .S0(n512), .Y(\normal/sll_15/n21 ) );
  MXI2X1 \normal/sll_15/U26  ( .A(\normal/sll_15/n22 ), .B(\normal/sll_15/n21 ), .S0(n503), .Y(\normal/N69 ) );
  MXI2X1 \normal/sll_15/U76  ( .A(\normal/sll_15/n65 ), .B(\normal/sll_15/n61 ), .S0(n512), .Y(\normal/sll_15/n18 ) );
  MXI2X1 \normal/sll_15/U29  ( .A(\normal/sll_15/n18 ), .B(\normal/sll_15/n17 ), .S0(n503), .Y(\normal/N66 ) );
  MXI2X1 \normal/sll_15/U28  ( .A(\normal/sll_15/n19 ), .B(\normal/sll_15/n18 ), .S0(n503), .Y(\normal/N67 ) );
  OAI21X1 \ctrl/add_1_root_add_16_2/U46  ( .A0(\ctrl/add_1_root_add_16_2/n49 ), 
        .A1(\ctrl/add_1_root_add_16_2/n41 ), .B0(
        \ctrl/add_1_root_add_16_2/n44 ), .Y(\ctrl/add_1_root_add_16_2/n40 ) );
  XOR2X1 \round/r298/U119  ( .A(\round/r298/n104 ), .B(\round/r298/n103 ), .Y(
        \round/N13 ) );
  XOR2X1 \round/r298/U68  ( .A(\round/r298/n62 ), .B(\round/r298/n61 ), .Y(
        \round/N21 ) );
  XOR2X1 \round/r298/U74  ( .A(\round/r298/n69 ), .B(\round/r298/n68 ), .Y(
        \round/N20 ) );
  XOR2X1 \round/r298/U82  ( .A(\round/r298/n74 ), .B(\round/r298/n73 ), .Y(
        \round/N19 ) );
  XNOR2X1 \round/r298/U96  ( .A(\round/r298/n84 ), .B(\round/r298/n83 ), .Y(
        \round/N17 ) );
  XOR2X1 \round/r298/U139  ( .A(\round/r298/n117 ), .B(n522), .Y(\round/N9 )
         );
  AO21X2 \mul/mult_6/U842  ( .A0(n700), .A1(sig_B[22]), .B0(n681), .Y(
        \mul/mult_6/n544 ) );
  AO21X2 \mul/mult_6/U759  ( .A0(n699), .A1(sig_B[22]), .B0(n683), .Y(
        \mul/mult_6/n540 ) );
  AOI21X1 \mul/mult_6/U754  ( .A0(\mul/mult_6/n30 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n539 ), .Y(\mul/mult_6/n1234 ) );
  AOI222XL \mul/mult_6/U380  ( .A0(n695), .A1(sig_B[11]), .B0(n696), .B1(
        sig_B[10]), .C0(\mul/mult_6/n78 ), .C1(sig_B[9]), .Y(\mul/mult_6/n987 ) );
  AOI21X1 \mul/mult_6/U675  ( .A0(\mul/mult_6/n40 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n536 ), .Y(\mul/mult_6/n1183 ) );
  OAI21X1 \mul/mult_6/U447  ( .A0(n570), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1034 ), .Y(\mul/mult_6/n1008 ) );
  XOR2X1 \mul/mult_6/U446  ( .A(\mul/mult_6/n1008 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n768 ) );
  AOI21X1 \mul/mult_6/U671  ( .A0(\mul/mult_6/n40 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n535 ), .Y(\mul/mult_6/n1182 ) );
  AO21X2 \mul/mult_6/U593  ( .A0(n518), .A1(sig_B[22]), .B0(n687), .Y(
        \mul/mult_6/n532 ) );
  AOI21X1 \mul/mult_6/U592  ( .A0(\mul/mult_6/n50 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n532 ), .Y(\mul/mult_6/n1131 ) );
  AOI21X1 \mul/mult_6/U588  ( .A0(\mul/mult_6/n50 ), .A1(sig_B[22]), .B0(n518), 
        .Y(\mul/mult_6/n1130 ) );
  AOI222XL \mul/mult_6/U362  ( .A0(n695), .A1(sig_B[17]), .B0(\mul/mult_6/n74 ), .B1(sig_B[16]), .C0(\mul/mult_6/n78 ), .C1(sig_B[15]), .Y(\mul/mult_6/n981 )
         );
  AO21X2 \mul/mult_6/U510  ( .A0(n690), .A1(sig_B[22]), .B0(n689), .Y(
        \mul/mult_6/n528 ) );
  AOI21X1 \mul/mult_6/U509  ( .A0(\mul/mult_6/n60 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n528 ), .Y(\mul/mult_6/n1079 ) );
  AOI21X1 \mul/mult_6/U426  ( .A0(\mul/mult_6/n70 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n524 ), .Y(\mul/mult_6/n1027 ) );
  AOI222XL \mul/mult_6/U350  ( .A0(\mul/mult_6/n72 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n74 ), .B1(sig_B[20]), .C0(\mul/mult_6/n78 ), .C1(
        sig_B[19]), .Y(\mul/mult_6/n977 ) );
  AOI222XL \mul/mult_6/U347  ( .A0(\mul/mult_6/n72 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n74 ), .B1(sig_B[21]), .C0(\mul/mult_6/n78 ), .C1(
        sig_B[20]), .Y(\mul/mult_6/n976 ) );
  AOI21X1 \mul/mult_6/U343  ( .A0(\mul/mult_6/n78 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n520 ), .Y(\mul/mult_6/n975 ) );
  OAI21X1 \mul/mult_6/U536  ( .A0(n571), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1088 ), .Y(\mul/mult_6/n1062 ) );
  XOR2X1 \mul/mult_6/U535  ( .A(\mul/mult_6/n1062 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n797 ) );
  OAI21X1 \mul/mult_6/U684  ( .A0(n591), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1186 ), .Y(\mul/mult_6/n1160 ) );
  XOR2X1 \mul/mult_6/U749  ( .A(\mul/mult_6/n1207 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n867 ) );
  XOR2X1 \mul/mult_6/U606  ( .A(\mul/mult_6/n1110 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n820 ) );
  OAI21X1 \mul/mult_6/U530  ( .A0(n570), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1086 ), .Y(\mul/mult_6/n1060 ) );
  XOR2X1 \mul/mult_6/U529  ( .A(\mul/mult_6/n1060 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n795 ) );
  XOR2X1 \mul/mult_6/U532  ( .A(\mul/mult_6/n1061 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n796 ) );
  XOR2X1 \mul/mult_6/U603  ( .A(\mul/mult_6/n1109 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n819 ) );
  OAI21X1 \mul/mult_6/U453  ( .A0(n571), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1036 ), .Y(\mul/mult_6/n1010 ) );
  XOR2X1 \mul/mult_6/U452  ( .A(\mul/mult_6/n1010 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n770 ) );
  XOR2X1 \mul/mult_6/U455  ( .A(\mul/mult_6/n1011 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n771 ) );
  OAI21X1 \mul/mult_6/U753  ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1234 ), .Y(\mul/mult_6/n1208 ) );
  XOR2X1 \mul/mult_6/U752  ( .A(\mul/mult_6/n1208 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n868 ) );
  OAI21X1 \mul/mult_6/U527  ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1085 ), .Y(\mul/mult_6/n1059 ) );
  XOR2X1 \mul/mult_6/U526  ( .A(\mul/mult_6/n1059 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n794 ) );
  XOR2X1 \mul/mult_6/U600  ( .A(\mul/mult_6/n1108 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n818 ) );
  XOR2X1 \mul/mult_6/U666  ( .A(\mul/mult_6/n1155 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n840 ) );
  XOR2X1 \mul/mult_6/U523  ( .A(\mul/mult_6/n1058 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n793 ) );
  OAI21X1 \mul/mult_6/U450  ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1035 ), .Y(\mul/mult_6/n1009 ) );
  XOR2X1 \mul/mult_6/U669  ( .A(\mul/mult_6/n1156 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n841 ) );
  XOR2X1 \mul/mult_6/U597  ( .A(\mul/mult_6/n1107 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n817 ) );
  OAI21X1 \mul/mult_6/U518  ( .A0(n591), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1082 ), .Y(\mul/mult_6/n1056 ) );
  XOR2X1 \mul/mult_6/U517  ( .A(\mul/mult_6/n1056 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n791 ) );
  XOR2X1 \mul/mult_6/U594  ( .A(\mul/mult_6/n1106 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n816 ) );
  XOR2X1 \mul/mult_6/U520  ( .A(\mul/mult_6/n1057 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n792 ) );
  XOR2X1 \mul/mult_6/U443  ( .A(\mul/mult_6/n1007 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n767 ) );
  OAI21X1 \mul/mult_6/U441  ( .A0(n569), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1032 ), .Y(\mul/mult_6/n1006 ) );
  XOR2X1 \mul/mult_6/U431  ( .A(\mul/mult_6/n1003 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n763 ) );
  NAND2X2 \expadd/add_0_root_sub_0_root_sub_8/U14  ( .A(
        \expadd/add_0_root_sub_0_root_sub_8/B[0] ), .B(exp_B[0]), .Y(
        \expadd/add_0_root_sub_0_root_sub_8/n11 ) );
  NAND2X2 \expadd/add_0_root_sub_0_root_sub_8/U11  ( .A(n657), .B(
        \expadd/add_0_root_sub_0_root_sub_8/n11 ), .Y(
        \expadd/add_0_root_sub_0_root_sub_8/n2 ) );
  NOR2BX8 \mul/mult_6/U1097  ( .AN(\mul/mult_6/n1443 ), .B(\mul/mult_6/n1451 ), 
        .Y(\mul/mult_6/n547 ) );
  ADDHX1 \selc/r299/U49  ( .A(\selc/r299/A[1] ), .B(\mul/mult_6/n125 ), .CO(
        \selc/r299/n48 ), .S(\selc/N114 ) );
  NAND2X2 \mul/mult_6/U1277  ( .A(sig_B[4]), .B(sig_B[5]), .Y(
        \mul/mult_6/n692 ) );
  NAND2X2 \mul/mult_6/U1228  ( .A(sig_B[10]), .B(sig_B[11]), .Y(
        \mul/mult_6/n661 ) );
  NAND2X2 \mul/mult_6/U1206  ( .A(sig_B[12]), .B(sig_B[13]), .Y(
        \mul/mult_6/n645 ) );
  NAND2X2 \mul/mult_6/U1165  ( .A(sig_B[16]), .B(sig_B[17]), .Y(
        \mul/mult_6/n616 ) );
  NAND2X2 \mul/mult_6/U1297  ( .A(\mul/mult_6/n731 ), .B(\mul/mult_6/n706 ), 
        .Y(\mul/mult_6/n572 ) );
  NOR2BX8 \mul/mult_6/U1083  ( .AN(\mul/mult_6/n1441 ), .B(\mul/mult_6/n1449 ), 
        .Y(\mul/mult_6/n539 ) );
  NAND2X2 \mul/mult_6/U1249  ( .A(\mul/mult_6/n725 ), .B(\mul/mult_6/n676 ), 
        .Y(\mul/mult_6/n566 ) );
  NAND2X2 \mul/mult_6/U1274  ( .A(\mul/mult_6/n728 ), .B(\mul/mult_6/n692 ), 
        .Y(\mul/mult_6/n569 ) );
  NOR2BX8 \mul/mult_6/U1090  ( .AN(\mul/mult_6/n1442 ), .B(\mul/mult_6/n1450 ), 
        .Y(\mul/mult_6/n543 ) );
  NAND2X2 \mul/mult_6/U1282  ( .A(\mul/mult_6/n729 ), .B(\mul/mult_6/n697 ), 
        .Y(\mul/mult_6/n570 ) );
  NAND2X2 \mul/mult_6/U1291  ( .A(\mul/mult_6/n730 ), .B(\mul/mult_6/n703 ), 
        .Y(\mul/mult_6/n571 ) );
  NAND2X2 \mul/mult_6/U1260  ( .A(\mul/mult_6/n726 ), .B(\mul/mult_6/n684 ), 
        .Y(\mul/mult_6/n567 ) );
  NAND2X2 \mul/mult_6/U1266  ( .A(\mul/mult_6/n727 ), .B(\mul/mult_6/n687 ), 
        .Y(\mul/mult_6/n568 ) );
  ADDHX1 \selc/r299/U48  ( .A(\selc/r299/A[2] ), .B(\selc/r299/n48 ), .CO(
        \selc/r299/n47 ), .S(\selc/N115 ) );
  ADDHX1 \selc/r299/U47  ( .A(\selc/r299/n47 ), .B(\selc/r299/A[3] ), .CO(
        \selc/r299/n46 ), .S(\selc/N116 ) );
  ADDHX1 \selc/r299/U46  ( .A(\selc/r299/n46 ), .B(\selc/r299/A[4] ), .CO(
        \selc/r299/n45 ), .S(\selc/N117 ) );
  ADDHX1 \selc/r299/U45  ( .A(\selc/r299/n45 ), .B(\selc/r299/A[5] ), .CO(
        \selc/r299/n44 ), .S(\selc/N118 ) );
  ADDHX1 \selc/r299/U44  ( .A(\selc/r299/n44 ), .B(\selc/r299/A[6] ), .CO(
        \selc/r299/n43 ), .S(\selc/N119 ) );
  ADDHX1 \selc/r299/U43  ( .A(\selc/r299/n43 ), .B(\selc/r299/A[7] ), .CO(
        \selc/r299/n42 ), .S(\selc/N120 ) );
  ADDHX1 \selc/r299/U42  ( .A(\selc/r299/n42 ), .B(\selc/r299/A[8] ), .CO(
        \selc/r299/n41 ), .S(\selc/N121 ) );
  ADDHX1 \selc/r299/U41  ( .A(\selc/r299/n41 ), .B(\selc/r299/A[9] ), .CO(
        \selc/r299/n40 ), .S(\selc/N122 ) );
  ADDHX1 \selc/r299/U40  ( .A(\selc/r299/n40 ), .B(\selc/r299/A[10] ), .CO(
        \selc/r299/n39 ), .S(\selc/N123 ) );
  ADDHX1 \selc/r299/U39  ( .A(\selc/r299/n39 ), .B(\selc/r299/A[11] ), .CO(
        \selc/r299/n38 ), .S(\selc/N124 ) );
  ADDHX1 \selc/r299/U38  ( .A(\selc/r299/n38 ), .B(\selc/r299/A[12] ), .CO(
        \selc/r299/n37 ), .S(\selc/N125 ) );
  ADDHX1 \selc/r299/U37  ( .A(\selc/r299/n37 ), .B(\selc/r299/A[13] ), .CO(
        \selc/r299/n36 ), .S(\selc/N126 ) );
  ADDHX1 \selc/r299/U36  ( .A(\selc/r299/n36 ), .B(\selc/r299/A[14] ), .CO(
        \selc/r299/n35 ), .S(\selc/N127 ) );
  ADDHX1 \selc/r299/U35  ( .A(\selc/r299/n35 ), .B(\selc/r299/A[15] ), .CO(
        \selc/r299/n34 ), .S(\selc/N128 ) );
  ADDHX1 \selc/r299/U34  ( .A(\selc/r299/n34 ), .B(\selc/r299/A[16] ), .CO(
        \selc/r299/n33 ), .S(\selc/N129 ) );
  ADDHX1 \selc/r299/U33  ( .A(\selc/r299/n33 ), .B(\selc/r299/A[17] ), .CO(
        \selc/r299/n32 ), .S(\selc/N130 ) );
  ADDHX1 \selc/r299/U32  ( .A(\selc/r299/n32 ), .B(\selc/r299/A[18] ), .CO(
        \selc/r299/n31 ), .S(\selc/N131 ) );
  ADDHX1 \selc/r299/U31  ( .A(\selc/r299/n31 ), .B(\selc/r299/A[19] ), .CO(
        \selc/r299/n30 ), .S(\selc/N132 ) );
  ADDHX1 \selc/r299/U30  ( .A(\selc/r299/n30 ), .B(\selc/r299/A[20] ), .CO(
        \selc/r299/n29 ), .S(\selc/N133 ) );
  ADDHX1 \selc/r299/U29  ( .A(\selc/r299/n29 ), .B(\selc/r299/A[21] ), .CO(
        \selc/r299/n28 ), .S(\selc/N134 ) );
  ADDHX1 \selc/r299/U28  ( .A(\selc/r299/n28 ), .B(\selc/r299/A[22] ), .CO(
        \selc/r299/n27 ), .S(\selc/N135 ) );
  ADDHX1 \selc/r299/U27  ( .A(\selc/r299/n27 ), .B(\selc/r299/A[23] ), .CO(
        \selc/r299/n26 ), .S(\selc/N136 ) );
  ADDHX1 \selc/r299/U26  ( .A(\selc/r299/n26 ), .B(\selc/r299/A[24] ), .CO(
        \selc/r299/n25 ), .S(\selc/N137 ) );
  ADDHX1 \selc/r299/U25  ( .A(\selc/r299/n25 ), .B(\selc/r299/A[25] ), .CO(
        \selc/r299/n24 ), .S(\selc/N138 ) );
  ADDHX1 \selc/r299/U24  ( .A(\selc/r299/n24 ), .B(\selc/r299/A[26] ), .CO(
        \selc/r299/n23 ), .S(\selc/N139 ) );
  ADDHX1 \selc/r299/U23  ( .A(\selc/r299/n23 ), .B(\selc/r299/A[27] ), .CO(
        \selc/r299/n22 ), .S(\selc/N140 ) );
  ADDHX1 \selc/r299/U22  ( .A(\selc/r299/n22 ), .B(\selc/r299/A[28] ), .CO(
        \selc/r299/n21 ), .S(\selc/N141 ) );
  ADDHX1 \selc/r299/U21  ( .A(\selc/r299/n21 ), .B(\selc/r299/A[29] ), .CO(
        \selc/r299/n20 ), .S(\selc/N142 ) );
  ADDHX1 \selc/r299/U20  ( .A(\selc/r299/n20 ), .B(\selc/r299/A[30] ), .CO(
        \selc/r299/n19 ), .S(\selc/N143 ) );
  ADDHX1 \selc/r299/U19  ( .A(\selc/r299/n19 ), .B(\selc/r299/A[31] ), .CO(
        \selc/r299/n18 ), .S(\selc/N144 ) );
  ADDHX1 \selc/r299/U18  ( .A(\selc/r299/n18 ), .B(\selc/r299/A[32] ), .CO(
        \selc/r299/n17 ), .S(\selc/N145 ) );
  ADDHX1 \selc/r299/U17  ( .A(\selc/r299/n17 ), .B(\selc/r299/A[33] ), .CO(
        \selc/r299/n16 ), .S(\selc/N146 ) );
  ADDHX1 \selc/r299/U16  ( .A(\selc/r299/n16 ), .B(\selc/r299/A[34] ), .CO(
        \selc/r299/n15 ), .S(\selc/N147 ) );
  ADDHX1 \selc/r299/U15  ( .A(\selc/r299/n15 ), .B(\selc/r299/A[35] ), .CO(
        \selc/r299/n14 ), .S(\selc/N148 ) );
  ADDHX1 \selc/r299/U14  ( .A(\selc/r299/n14 ), .B(\selc/r299/A[36] ), .CO(
        \selc/r299/n13 ), .S(\selc/N149 ) );
  ADDHX1 \selc/r299/U13  ( .A(\selc/r299/n13 ), .B(\selc/r299/A[37] ), .CO(
        \selc/r299/n12 ), .S(\selc/N150 ) );
  ADDHX1 \selc/r299/U12  ( .A(\selc/r299/n12 ), .B(\selc/r299/A[38] ), .CO(
        \selc/r299/n11 ), .S(\selc/N151 ) );
  ADDHX1 \selc/r299/U11  ( .A(\selc/r299/n11 ), .B(\selc/r299/A[39] ), .CO(
        \selc/r299/n10 ), .S(\selc/N152 ) );
  ADDHX1 \selc/r299/U10  ( .A(\selc/r299/n10 ), .B(\selc/r299/A[40] ), .CO(
        \selc/r299/n9 ), .S(\selc/N153 ) );
  ADDHX1 \selc/r300/U1_1_24  ( .A(\selc/r300/A[24] ), .B(\selc/r300/carry[24] ), .CO(\selc/r300/carry[25] ), .S(\selc/N187 ) );
  ADDHX1 \selc/r300/U1_1_25  ( .A(\selc/r300/A[25] ), .B(\selc/r300/carry[25] ), .CO(\selc/r300/carry[26] ), .S(\selc/N188 ) );
  ADDHX1 \selc/r300/U1_1_26  ( .A(\selc/r300/A[26] ), .B(\selc/r300/carry[26] ), .CO(\selc/r300/carry[27] ), .S(\selc/N189 ) );
  ADDHX1 \selc/r300/U1_1_27  ( .A(\selc/r300/A[27] ), .B(\selc/r300/carry[27] ), .CO(\selc/r300/carry[28] ), .S(\selc/N190 ) );
  ADDHX1 \selc/r300/U1_1_28  ( .A(\selc/r300/A[28] ), .B(\selc/r300/carry[28] ), .CO(\selc/r300/carry[29] ), .S(\selc/N191 ) );
  ADDHX1 \selc/r300/U1_1_29  ( .A(\selc/r300/A[29] ), .B(\selc/r300/carry[29] ), .CO(\selc/r300/carry[30] ), .S(\selc/N192 ) );
  ADDHX1 \selc/r300/U1_1_30  ( .A(\selc/r300/A[30] ), .B(\selc/r300/carry[30] ), .CO(\selc/r300/carry[31] ), .S(\selc/N193 ) );
  ADDHX1 \selc/r300/U1_1_31  ( .A(\selc/r300/A[31] ), .B(\selc/r300/carry[31] ), .CO(\selc/r300/carry[32] ), .S(\selc/N194 ) );
  ADDHX1 \selc/r300/U1_1_32  ( .A(\selc/r300/A[32] ), .B(\selc/r300/carry[32] ), .CO(\selc/r300/carry[33] ), .S(\selc/N195 ) );
  ADDHX1 \selc/r300/U1_1_33  ( .A(\selc/r300/A[33] ), .B(\selc/r300/carry[33] ), .CO(\selc/r300/carry[34] ), .S(\selc/N196 ) );
  ADDHX1 \selc/r300/U1_1_34  ( .A(\selc/r300/A[34] ), .B(\selc/r300/carry[34] ), .CO(\selc/r300/carry[35] ), .S(\selc/N197 ) );
  ADDHX1 \selc/r300/U1_1_35  ( .A(\selc/r300/A[35] ), .B(\selc/r300/carry[35] ), .CO(\selc/r300/carry[36] ), .S(\selc/N198 ) );
  ADDHX1 \selc/r300/U1_1_36  ( .A(\selc/r300/A[36] ), .B(\selc/r300/carry[36] ), .CO(\selc/r300/carry[37] ), .S(\selc/N199 ) );
  ADDHX1 \selc/r300/U1_1_37  ( .A(\selc/r300/A[37] ), .B(\selc/r300/carry[37] ), .CO(\selc/r300/carry[38] ), .S(\selc/N200 ) );
  ADDHX1 \selc/r300/U1_1_38  ( .A(\selc/r300/A[38] ), .B(\selc/r300/carry[38] ), .CO(\selc/r300/carry[39] ), .S(\selc/N201 ) );
  ADDHX1 \selc/r300/U1_1_39  ( .A(\selc/r300/A[39] ), .B(\selc/r300/carry[39] ), .CO(\selc/r300/carry[40] ), .S(\selc/N202 ) );
  ADDHX1 \selc/r300/U1_1_40  ( .A(\selc/r300/A[40] ), .B(\selc/r300/carry[40] ), .CO(\selc/r300/carry[41] ), .S(\selc/N203 ) );
  ADDHX1 \selc/r300/U1_1_41  ( .A(\selc/r300/A[41] ), .B(\selc/r300/carry[41] ), .CO(\selc/r300/carry[42] ), .S(\selc/N204 ) );
  ADDHX1 \selc/r300/U1_1_42  ( .A(\selc/r300/A[42] ), .B(\selc/r300/carry[42] ), .CO(\selc/r300/carry[43] ), .S(\selc/N205 ) );
  ADDHX1 \selc/r300/U1_1_43  ( .A(\selc/r300/A[43] ), .B(\selc/r300/carry[43] ), .CO(\selc/r300/carry[44] ), .S(\selc/N206 ) );
  ADDHX1 \selc/r300/U1_1_44  ( .A(\selc/r300/A[44] ), .B(\selc/r300/carry[44] ), .CO(\selc/r300/carry[45] ), .S(\selc/N207 ) );
  ADDHX1 \selc/r300/U1_1_45  ( .A(\selc/r300/A[45] ), .B(\selc/r300/carry[45] ), .CO(\selc/N209 ), .S(\selc/N208 ) );
  NOR2X2 \sigadd/add_9/U340  ( .A(ali_P[1]), .B(ali_C[1]), .Y(
        \sigadd/add_9/n243 ) );
  NAND2X2 \sigadd/add_9/U341  ( .A(ali_P[1]), .B(ali_C[1]), .Y(
        \sigadd/add_9/n244 ) );
  NAND2X2 \sigadd/add_9/U335  ( .A(ali_P[2]), .B(ali_C[2]), .Y(
        \sigadd/add_9/n241 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U49  ( .A(\sigadd/add_9/n50 ), .B(
        \sigadd/sub_add_11_b0/n98 ), .CO(\sigadd/sub_add_11_b0/n48 ), .S(
        \sigadd/N3 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U48  ( .A(\sigadd/sub_add_11_b0/n97 ), .B(
        \sigadd/sub_add_11_b0/n48 ), .CO(\sigadd/sub_add_11_b0/n47 ), .S(
        \sigadd/N4 ) );
  NOR2X2 \sigadd/add_9/U326  ( .A(ali_P[3]), .B(ali_C[3]), .Y(
        \sigadd/add_9/n235 ) );
  NAND2X2 \sigadd/add_9/U327  ( .A(ali_P[3]), .B(ali_C[3]), .Y(
        \sigadd/add_9/n236 ) );
  NAND2X2 \sigadd/add_9/U321  ( .A(ali_P[4]), .B(ali_C[4]), .Y(
        \sigadd/add_9/n233 ) );
  NOR2X2 \sigadd/add_9/U312  ( .A(ali_P[5]), .B(ali_C[5]), .Y(
        \sigadd/add_9/n227 ) );
  NAND2X2 \sigadd/add_9/U313  ( .A(ali_P[5]), .B(ali_C[5]), .Y(
        \sigadd/add_9/n228 ) );
  NAND2X2 \sigadd/add_9/U307  ( .A(ali_P[6]), .B(ali_C[6]), .Y(
        \sigadd/add_9/n225 ) );
  NOR2X2 \sigadd/add_9/U298  ( .A(ali_P[7]), .B(ali_C[7]), .Y(
        \sigadd/add_9/n219 ) );
  NAND2X2 \sigadd/add_9/U299  ( .A(ali_P[7]), .B(ali_C[7]), .Y(
        \sigadd/add_9/n220 ) );
  NAND2X2 \sigadd/add_9/U293  ( .A(ali_P[8]), .B(ali_C[8]), .Y(
        \sigadd/add_9/n217 ) );
  NOR2X2 \sigadd/add_9/U284  ( .A(ali_P[9]), .B(ali_C[9]), .Y(
        \sigadd/add_9/n211 ) );
  NAND2X2 \sigadd/add_9/U285  ( .A(ali_P[9]), .B(ali_C[9]), .Y(
        \sigadd/add_9/n212 ) );
  NAND2X2 \sigadd/add_9/U279  ( .A(ali_P[10]), .B(ali_C[10]), .Y(
        \sigadd/add_9/n209 ) );
  NAND2X2 \sigadd/add_9/U271  ( .A(ali_P[11]), .B(ali_C[11]), .Y(
        \sigadd/add_9/n204 ) );
  NAND2X2 \sigadd/add_9/U265  ( .A(ali_P[12]), .B(ali_C[12]), .Y(
        \sigadd/add_9/n201 ) );
  NAND2X2 \sigadd/add_9/U125  ( .A(ali_P[32]), .B(ali_C[32]), .Y(
        \sigadd/add_9/n121 ) );
  NAND2X2 \sigadd/add_9/U111  ( .A(ali_P[34]), .B(ali_C[34]), .Y(
        \sigadd/add_9/n113 ) );
  NAND2X2 \sigadd/add_9/U97  ( .A(ali_P[36]), .B(ali_C[36]), .Y(
        \sigadd/add_9/n105 ) );
  NAND2X2 \sigadd/add_9/U83  ( .A(ali_P[38]), .B(ali_C[38]), .Y(
        \sigadd/add_9/n97 ) );
  NAND2X2 \sigadd/add_9/U69  ( .A(ali_P[40]), .B(ali_C[40]), .Y(
        \sigadd/add_9/n89 ) );
  NAND2X2 \sigadd/add_9/U55  ( .A(ali_P[42]), .B(ali_C[42]), .Y(
        \sigadd/add_9/n81 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U47  ( .A(\sigadd/sub_add_11_b0/n96 ), .B(
        \sigadd/sub_add_11_b0/n47 ), .CO(\sigadd/sub_add_11_b0/n46 ), .S(
        \sigadd/N5 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U46  ( .A(\sigadd/sub_add_11_b0/n95 ), .B(
        \sigadd/sub_add_11_b0/n46 ), .CO(\sigadd/sub_add_11_b0/n45 ), .S(
        \sigadd/N6 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U45  ( .A(n656), .B(\sigadd/sub_add_11_b0/n45 ), 
        .CO(\sigadd/sub_add_11_b0/n44 ), .S(\sigadd/N7 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U44  ( .A(n649), .B(\sigadd/sub_add_11_b0/n44 ), 
        .CO(\sigadd/sub_add_11_b0/n43 ), .S(\sigadd/N8 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U43  ( .A(n648), .B(\sigadd/sub_add_11_b0/n43 ), 
        .CO(\sigadd/sub_add_11_b0/n42 ), .S(\sigadd/N9 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U42  ( .A(n636), .B(\sigadd/sub_add_11_b0/n42 ), 
        .CO(\sigadd/sub_add_11_b0/n41 ), .S(\sigadd/N10 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U41  ( .A(n647), .B(\sigadd/sub_add_11_b0/n41 ), 
        .CO(\sigadd/sub_add_11_b0/n40 ), .S(\sigadd/N11 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U40  ( .A(n635), .B(\sigadd/sub_add_11_b0/n40 ), 
        .CO(\sigadd/sub_add_11_b0/n39 ), .S(\sigadd/N12 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U36  ( .A(n633), .B(\sigadd/sub_add_11_b0/n36 ), 
        .CO(\sigadd/sub_add_11_b0/n35 ), .S(\sigadd/N16 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U35  ( .A(n644), .B(\sigadd/sub_add_11_b0/n35 ), 
        .CO(\sigadd/sub_add_11_b0/n34 ), .S(\sigadd/N17 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U34  ( .A(n623), .B(\sigadd/sub_add_11_b0/n34 ), 
        .CO(\sigadd/sub_add_11_b0/n33 ), .S(\sigadd/N18 ) );
  ADDHX1 \sigadd/sub_add_11_b0/U27  ( .A(n616), .B(\sigadd/sub_add_11_b0/n27 ), 
        .CO(\sigadd/sub_add_11_b0/n26 ), .S(\sigadd/N25 ) );
  NAND2BX2 \normal/srl_15/U257  ( .AN(n703), .B(add_out[37]), .Y(
        \normal/srl_15/n236 ) );
  NAND2BX2 \normal/srl_15/U255  ( .AN(n703), .B(add_out[39]), .Y(
        \normal/srl_15/n238 ) );
  NAND2BX2 \normal/srl_15/U157  ( .AN(n504), .B(\normal/srl_15/n186 ), .Y(
        \normal/srl_15/n136 ) );
  NAND2BX2 \normal/srl_15/U249  ( .AN(n703), .B(add_out[45]), .Y(
        \normal/srl_15/n244 ) );
  NAND2BX2 \normal/srl_15/U247  ( .AN(n703), .B(add_out[47]), .Y(
        \normal/srl_15/n246 ) );
  NAND2BX2 \normal/srl_15/U149  ( .AN(n504), .B(\normal/srl_15/n194 ), .Y(
        \normal/srl_15/n144 ) );
  NAND2BX2 \normal/srl_15/U253  ( .AN(n703), .B(\normal/srl_15/A[41] ), .Y(
        \normal/srl_15/n240 ) );
  NAND2BX2 \normal/srl_15/U251  ( .AN(n703), .B(add_out[43]), .Y(
        \normal/srl_15/n242 ) );
  NAND2BX2 \normal/srl_15/U153  ( .AN(n504), .B(\normal/srl_15/n190 ), .Y(
        \normal/srl_15/n140 ) );
  NAND2BX2 \normal/srl_15/U245  ( .AN(n703), .B(add_out[49]), .Y(
        \normal/srl_15/n248 ) );
  NOR2X2 \normal/srl_15/U195  ( .A(n514), .B(\normal/srl_15/n248 ), .Y(
        \normal/srl_15/n198 ) );
  NAND2BX2 \normal/srl_15/U145  ( .AN(n504), .B(\normal/srl_15/n198 ), .Y(
        \normal/srl_15/n148 ) );
  NAND2BX2 \normal/srl_15/U256  ( .AN(n703), .B(add_out[38]), .Y(
        \normal/srl_15/n237 ) );
  NAND2BX2 \normal/srl_15/U254  ( .AN(n703), .B(\normal/srl_15/A[40] ), .Y(
        \normal/srl_15/n239 ) );
  NAND2BX2 \normal/srl_15/U156  ( .AN(n504), .B(\normal/srl_15/n187 ), .Y(
        \normal/srl_15/n137 ) );
  NAND2BX2 \normal/srl_15/U248  ( .AN(n703), .B(add_out[46]), .Y(
        \normal/srl_15/n245 ) );
  NAND2BX2 \normal/srl_15/U148  ( .AN(n504), .B(\normal/srl_15/n195 ), .Y(
        \normal/srl_15/n145 ) );
  NAND2BX2 \normal/srl_15/U252  ( .AN(n703), .B(add_out[42]), .Y(
        \normal/srl_15/n241 ) );
  NAND2BX2 \normal/srl_15/U250  ( .AN(n703), .B(\normal/srl_15/A[44] ), .Y(
        \normal/srl_15/n243 ) );
  NAND2BX2 \normal/srl_15/U152  ( .AN(n504), .B(\normal/srl_15/n191 ), .Y(
        \normal/srl_15/n141 ) );
  NOR2X2 \normal/srl_15/U102  ( .A(\normal/srl_15/n141 ), .B(n513), .Y(
        \normal/srl_15/n91 ) );
  NAND2BX2 \normal/sll_15/U276  ( .AN(n714), .B(add_out[5]), .Y(
        \normal/sll_15/n194 ) );
  NAND2BX2 \normal/sll_15/U278  ( .AN(n714), .B(add_out[3]), .Y(
        \normal/sll_15/n192 ) );
  NAND2BX2 \normal/sll_15/U280  ( .AN(n703), .B(\normal/srl_15/A[1] ), .Y(
        \normal/sll_15/n190 ) );
  NOR2X2 \normal/sll_15/U233  ( .A(n715), .B(\normal/sll_15/n190 ), .Y(
        \normal/sll_15/n143 ) );
  NAND2BX2 \normal/sll_15/U162  ( .AN(n504), .B(\normal/sll_15/n167 ), .Y(
        \normal/sll_15/n120 ) );
  NAND2BX2 \normal/sll_15/U277  ( .AN(n714), .B(\normal/srl_15/A[4] ), .Y(
        \normal/sll_15/n193 ) );
  NAND2BX2 \normal/sll_15/U279  ( .AN(n703), .B(add_out[2]), .Y(
        \normal/sll_15/n191 ) );
  NAND2BX2 \normal/sll_15/U159  ( .AN(n504), .B(\normal/sll_15/n170 ), .Y(
        \normal/sll_15/n123 ) );
  NAND2BX2 \normal/sll_15/U281  ( .AN(n703), .B(\sigadd/sig[0] ), .Y(
        \normal/sll_15/n189 ) );
  NOR2X2 \normal/sll_15/U234  ( .A(n715), .B(\normal/sll_15/n189 ), .Y(
        \normal/sll_15/n142 ) );
  NAND2BX2 \normal/srl_15/U258  ( .AN(n703), .B(\normal/srl_15/A[36] ), .Y(
        \normal/srl_15/n235 ) );
  NAND2BX2 \normal/srl_15/U158  ( .AN(n504), .B(\normal/srl_15/n185 ), .Y(
        \normal/srl_15/n135 ) );
  NAND2BX2 \normal/srl_15/U150  ( .AN(n504), .B(\normal/srl_15/n193 ), .Y(
        \normal/srl_15/n143 ) );
  NAND2BX2 \normal/srl_15/U154  ( .AN(n504), .B(\normal/srl_15/n189 ), .Y(
        \normal/srl_15/n139 ) );
  NOR2X2 \normal/srl_15/U196  ( .A(n514), .B(\normal/srl_15/n247 ), .Y(
        \normal/srl_15/n197 ) );
  NAND2BX2 \normal/srl_15/U146  ( .AN(n504), .B(\normal/srl_15/n197 ), .Y(
        \normal/srl_15/n147 ) );
  NAND2BX2 \normal/sll_15/U160  ( .AN(n504), .B(\normal/sll_15/n169 ), .Y(
        \normal/sll_15/n122 ) );
  NAND2BX2 \normal/sll_15/U156  ( .AN(n504), .B(\normal/sll_15/n173 ), .Y(
        \normal/sll_15/n126 ) );
  NAND2BX2 \normal/srl_15/U155  ( .AN(n504), .B(\normal/srl_15/n188 ), .Y(
        \normal/srl_15/n138 ) );
  NAND2BX2 \normal/srl_15/U147  ( .AN(n504), .B(\normal/srl_15/n196 ), .Y(
        \normal/srl_15/n146 ) );
  NAND2BX2 \normal/srl_15/U151  ( .AN(n504), .B(\normal/srl_15/n192 ), .Y(
        \normal/srl_15/n142 ) );
  NOR2X2 \normal/srl_15/U101  ( .A(\normal/srl_15/n142 ), .B(n513), .Y(
        \normal/srl_15/n92 ) );
  NAND2BX2 \normal/sll_15/U275  ( .AN(n714), .B(\normal/srl_15/A[6] ), .Y(
        \normal/sll_15/n195 ) );
  NAND2BX2 \normal/sll_15/U161  ( .AN(n504), .B(\normal/sll_15/n168 ), .Y(
        \normal/sll_15/n121 ) );
  NOR2X2 \normal/srl_15/U100  ( .A(\normal/srl_15/n143 ), .B(n513), .Y(
        \normal/srl_15/n93 ) );
  NAND2BX2 \normal/sll_15/U274  ( .AN(n714), .B(add_out[7]), .Y(
        \normal/sll_15/n196 ) );
  NAND2BX2 \normal/srl_15/U259  ( .AN(n703), .B(add_out[35]), .Y(
        \normal/srl_15/n234 ) );
  NAND2BX2 \normal/srl_15/U159  ( .AN(n504), .B(\normal/srl_15/n184 ), .Y(
        \normal/srl_15/n134 ) );
  NAND2BX2 \normal/srl_15/U260  ( .AN(n703), .B(add_out[34]), .Y(
        \normal/srl_15/n233 ) );
  NAND2BX2 \normal/srl_15/U160  ( .AN(n504), .B(\normal/srl_15/n183 ), .Y(
        \normal/srl_15/n133 ) );
  NAND2BX2 \normal/srl_15/U162  ( .AN(n504), .B(\normal/srl_15/n181 ), .Y(
        \normal/srl_15/n131 ) );
  NAND2BX2 \normal/srl_15/U161  ( .AN(n504), .B(\normal/srl_15/n182 ), .Y(
        \normal/srl_15/n132 ) );
  NAND2BX2 \normal/sll_15/U266  ( .AN(n714), .B(add_out[15]), .Y(
        \normal/sll_15/n204 ) );
  NAND2BX2 \normal/sll_15/U267  ( .AN(n714), .B(add_out[14]), .Y(
        \normal/sll_15/n203 ) );
  NAND2BX2 \normal/sll_15/U171  ( .AN(n504), .B(\normal/sll_15/n158 ), .Y(
        \normal/sll_15/n111 ) );
  NAND2BX2 \normal/sll_15/U268  ( .AN(n714), .B(add_out[13]), .Y(
        \normal/sll_15/n202 ) );
  NAND2BX2 \normal/sll_15/U172  ( .AN(n504), .B(\normal/sll_15/n157 ), .Y(
        \normal/sll_15/n110 ) );
  NAND2BX2 \normal/srl_15/U170  ( .AN(n504), .B(\normal/srl_15/n173 ), .Y(
        \normal/srl_15/n123 ) );
  NAND2BX2 \normal/sll_15/U270  ( .AN(n714), .B(\normal/srl_15/A[11] ), .Y(
        \normal/sll_15/n200 ) );
  NAND2BX2 \normal/sll_15/U272  ( .AN(n714), .B(\normal/srl_15/A[9] ), .Y(
        \normal/sll_15/n198 ) );
  NAND2BX2 \normal/sll_15/U176  ( .AN(n504), .B(\normal/sll_15/n153 ), .Y(
        \normal/sll_15/n106 ) );
  NAND2BX2 \normal/sll_15/U269  ( .AN(n714), .B(\normal/srl_15/A[12] ), .Y(
        \normal/sll_15/n201 ) );
  NAND2BX2 \normal/sll_15/U173  ( .AN(n504), .B(\normal/sll_15/n156 ), .Y(
        \normal/sll_15/n109 ) );
  NAND2BX2 \normal/sll_15/U271  ( .AN(n714), .B(\normal/srl_15/A[10] ), .Y(
        \normal/sll_15/n199 ) );
  NAND2BX2 \normal/sll_15/U273  ( .AN(n714), .B(\normal/srl_15/A[8] ), .Y(
        \normal/sll_15/n197 ) );
  NAND2BX2 \normal/sll_15/U177  ( .AN(n504), .B(\normal/sll_15/n152 ), .Y(
        \normal/sll_15/n105 ) );
  NAND2BX2 \normal/srl_15/U169  ( .AN(n504), .B(\normal/srl_15/n174 ), .Y(
        \normal/srl_15/n124 ) );
  NAND2BX2 \normal/sll_15/U175  ( .AN(n504), .B(\normal/sll_15/n154 ), .Y(
        \normal/sll_15/n107 ) );
  NAND2BX2 \normal/srl_15/U168  ( .AN(n504), .B(\normal/srl_15/n175 ), .Y(
        \normal/srl_15/n125 ) );
  NAND2BX2 \normal/sll_15/U174  ( .AN(n504), .B(\normal/sll_15/n155 ), .Y(
        \normal/sll_15/n108 ) );
  NOR2X2 \normal/srl_15/U99  ( .A(\normal/srl_15/n144 ), .B(n513), .Y(
        \normal/srl_15/n94 ) );
  NOR2X2 \normal/srl_15/U98  ( .A(\normal/srl_15/n145 ), .B(n513), .Y(
        \normal/srl_15/n95 ) );
  NAND2BX2 \normal/srl_15/U48  ( .AN(n704), .B(\normal/srl_15/n95 ), .Y(
        \normal/srl_15/n47 ) );
  NOR2X2 \normal/srl_15/U97  ( .A(\normal/srl_15/n146 ), .B(n513), .Y(
        \normal/srl_15/n96 ) );
  NAND2BX2 \normal/srl_15/U47  ( .AN(n704), .B(\normal/srl_15/n96 ), .Y(
        \normal/srl_15/n48 ) );
  NAND2BX2 \normal/srl_15/U174  ( .AN(n504), .B(\normal/srl_15/n169 ), .Y(
        \normal/srl_15/n119 ) );
  NAND2BX2 \normal/sll_15/U178  ( .AN(n504), .B(\normal/sll_15/n151 ), .Y(
        \normal/sll_15/n104 ) );
  NAND2BX2 \normal/sll_15/U186  ( .AN(n504), .B(\normal/sll_15/n143 ), .Y(
        \normal/sll_15/n96 ) );
  NAND2BX2 \normal/sll_15/U182  ( .AN(n504), .B(\normal/sll_15/n147 ), .Y(
        \normal/sll_15/n100 ) );
  NOR2X2 \normal/sll_15/U135  ( .A(\normal/sll_15/n100 ), .B(n513), .Y(
        \normal/sll_15/n53 ) );
  NAND2BX2 \normal/sll_15/U179  ( .AN(n504), .B(\normal/sll_15/n150 ), .Y(
        \normal/sll_15/n103 ) );
  NAND2BX2 \normal/sll_15/U187  ( .AN(n504), .B(\normal/sll_15/n142 ), .Y(
        \normal/sll_15/n95 ) );
  NAND2BX2 \normal/sll_15/U183  ( .AN(n504), .B(\normal/sll_15/n146 ), .Y(
        \normal/sll_15/n99 ) );
  NOR2X2 \normal/sll_15/U136  ( .A(\normal/sll_15/n99 ), .B(n513), .Y(
        \normal/sll_15/n52 ) );
  NAND2BX2 \normal/sll_15/U185  ( .AN(n504), .B(\normal/sll_15/n144 ), .Y(
        \normal/sll_15/n97 ) );
  NAND2BX2 \normal/sll_15/U181  ( .AN(n504), .B(\normal/sll_15/n148 ), .Y(
        \normal/sll_15/n101 ) );
  NOR2X2 \normal/sll_15/U134  ( .A(\normal/sll_15/n101 ), .B(n513), .Y(
        \normal/sll_15/n54 ) );
  NAND2BX2 \normal/sll_15/U184  ( .AN(n504), .B(\normal/sll_15/n145 ), .Y(
        \normal/sll_15/n98 ) );
  NAND2BX2 \normal/sll_15/U180  ( .AN(n504), .B(\normal/sll_15/n149 ), .Y(
        \normal/sll_15/n102 ) );
  NOR2X2 \normal/sll_15/U133  ( .A(\normal/sll_15/n102 ), .B(n513), .Y(
        \normal/sll_15/n55 ) );
  NOR2X2 \normal/sll_15/U139  ( .A(\normal/sll_15/n96 ), .B(n513), .Y(
        \normal/sll_15/n49 ) );
  NOR2X2 \normal/sll_15/U140  ( .A(\normal/sll_15/n95 ), .B(n513), .Y(
        \normal/sll_15/n48 ) );
  NOR2X2 \normal/sll_15/U138  ( .A(\normal/sll_15/n97 ), .B(n513), .Y(
        \normal/sll_15/n50 ) );
  NOR2X2 \normal/sll_15/U137  ( .A(\normal/sll_15/n98 ), .B(n513), .Y(
        \normal/sll_15/n51 ) );
  NAND2BX2 \normal/sll_15/U93  ( .AN(n704), .B(\normal/sll_15/n48 ), .Y(
        \normal/sll_15/n1 ) );
  NAND2X2 \ctrl/add_1_root_add_16_2/U23  ( .A(\ctrl/add_1_root_add_16_2/n30 ), 
        .B(n533), .Y(\ctrl/add_1_root_add_16_2/n23 ) );
  NAND2X2 \ctrl/add_1_root_add_16_2/U52  ( .A(n704), .B(
        \ctrl/add_1_root_add_16_2/A[2] ), .Y(\ctrl/add_1_root_add_16_2/n44 )
         );
  NAND2X2 \ctrl/add_1_root_add_16_2/U42  ( .A(n513), .B(mux_out[3]), .Y(
        \ctrl/add_1_root_add_16_2/n37 ) );
  NAND2X2 \ctrl/add_1_root_add_16_2/U30  ( .A(n703), .B(
        \ctrl/add_1_root_add_16_2/A[4] ), .Y(\ctrl/add_1_root_add_16_2/n28 )
         );
  NAND2X2 \ctrl/sub_0_root_add_0_root_sub_16/U29  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/n38 ), .B(
        \ctrl/sub_0_root_add_0_root_sub_16/n26 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n4 ) );
  NOR2X2 \ctrl/add_1_root_add_16_2/U45  ( .A(\ctrl/add_1_root_add_16_2/n48 ), 
        .B(\ctrl/add_1_root_add_16_2/n41 ), .Y(\ctrl/add_1_root_add_16_2/n39 )
         );
  NAND2X2 \ctrl/add_1_root_add_16_2/U39  ( .A(\ctrl/add_1_root_add_16_2/n67 ), 
        .B(\ctrl/add_1_root_add_16_2/n37 ), .Y(\ctrl/add_1_root_add_16_2/n3 )
         );
  NAND2X2 \ctrl/sub_0_root_add_0_root_sub_16/U43  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/n40 ), .B(
        \ctrl/sub_0_root_add_0_root_sub_16/n34 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n6 ) );
  NOR2X2 \round/r298/U56  ( .A(\round/r298/n47 ), .B(\round/r298/n64 ), .Y(
        \round/r298/n46 ) );
  NAND2X2 \round/r298/U55  ( .A(\round/r298/n46 ), .B(\round/r298/n84 ), .Y(
        \round/r298/n45 ) );
  NAND2X2 \round/r298/U61  ( .A(\round/r298/n51 ), .B(\round/r298/n84 ), .Y(
        \round/r298/n50 ) );
  NOR2X2 \round/r298/U70  ( .A(\round/r298/n64 ), .B(\round/r298/n61 ), .Y(
        \round/r298/n58 ) );
  NAND2X2 \round/r298/U69  ( .A(\round/r298/n58 ), .B(\round/r298/n84 ), .Y(
        \round/r298/n57 ) );
  NAND2X2 \round/r298/U83  ( .A(\round/r298/n84 ), .B(\round/r298/n70 ), .Y(
        \round/r298/n69 ) );
  NAND2X2 \round/r298/U89  ( .A(\round/r298/n84 ), .B(\round/r298/n75 ), .Y(
        \round/r298/n74 ) );
  NAND2X2 \round/r298/U97  ( .A(\round/r298/n84 ), .B(norm_out[12]), .Y(
        \round/r298/n81 ) );
  NOR2BX8 \mul/mult_6/U1076  ( .AN(\mul/mult_6/n1440 ), .B(\mul/mult_6/n1448 ), 
        .Y(\mul/mult_6/n535 ) );
  NAND2X2 \mul/mult_6/U1211  ( .A(\mul/mult_6/n721 ), .B(\mul/mult_6/n650 ), 
        .Y(\mul/mult_6/n562 ) );
  NAND2X2 \mul/mult_6/U1225  ( .A(\mul/mult_6/n722 ), .B(\mul/mult_6/n661 ), 
        .Y(\mul/mult_6/n563 ) );
  NOR2BX8 \mul/mult_6/U1062  ( .AN(\mul/mult_6/n1438 ), .B(\mul/mult_6/n1446 ), 
        .Y(\mul/mult_6/n54 ) );
  NAND2X2 \mul/mult_6/U1203  ( .A(\mul/mult_6/n720 ), .B(\mul/mult_6/n645 ), 
        .Y(\mul/mult_6/n561 ) );
  NAND2X2 \mul/mult_6/U1191  ( .A(\mul/mult_6/n719 ), .B(\mul/mult_6/n636 ), 
        .Y(\mul/mult_6/n560 ) );
  NOR2BX8 \mul/mult_6/U1055  ( .AN(\mul/mult_6/n1437 ), .B(\mul/mult_6/n1445 ), 
        .Y(\mul/mult_6/n64 ) );
  NAND2X2 \mul/mult_6/U1183  ( .A(\mul/mult_6/n718 ), .B(\mul/mult_6/n631 ), 
        .Y(\mul/mult_6/n559 ) );
  NAND2X2 \mul/mult_6/U1170  ( .A(\mul/mult_6/n717 ), .B(\mul/mult_6/n621 ), 
        .Y(\mul/mult_6/n558 ) );
  NAND2X2 \mul/mult_6/U1162  ( .A(\mul/mult_6/n716 ), .B(\mul/mult_6/n616 ), 
        .Y(\mul/mult_6/n557 ) );
  NAND2X2 \mul/mult_6/U1152  ( .A(\mul/mult_6/n715 ), .B(\mul/mult_6/n609 ), 
        .Y(\mul/mult_6/n556 ) );
  NAND2X2 \mul/mult_6/U1134  ( .A(\mul/mult_6/n713 ), .B(\mul/mult_6/n597 ), 
        .Y(\mul/mult_6/n554 ) );
  NAND2X2 \mul/mult_6/U1144  ( .A(\mul/mult_6/n714 ), .B(\mul/mult_6/n604 ), 
        .Y(\mul/mult_6/n555 ) );
  NAND2X2 \mul/mult_6/U1126  ( .A(\mul/mult_6/n712 ), .B(\mul/mult_6/n592 ), 
        .Y(\mul/mult_6/n553 ) );
  NAND2X2 \mul/mult_6/U1118  ( .A(n592), .B(\mul/mult_6/n587 ), .Y(
        \mul/mult_6/n552 ) );
  NOR2X8 \round/r298/U48  ( .A(\round/r298/n40 ), .B(\round/r298/n85 ), .Y(
        \round/r298/n1 ) );
  AOI222XL \mul/mult_6/U685  ( .A0(\mul/mult_6/n32 ), .A1(sig_B[20]), .B0(n698), .B1(sig_B[19]), .C0(\mul/mult_6/n40 ), .C1(sig_B[18]), .Y(\mul/mult_6/n1186 ) );
  XOR2X1 \mul/mult_6/U458  ( .A(\mul/mult_6/n1012 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n772 ) );
  AOI222XL \mul/mult_6/U679  ( .A0(\mul/mult_6/n32 ), .A1(sig_B[22]), .B0(n698), .B1(sig_B[21]), .C0(\mul/mult_6/n40 ), .C1(sig_B[20]), .Y(\mul/mult_6/n1184 ) );
  AOI222XL \mul/mult_6/U519  ( .A0(\mul/mult_6/n52 ), .A1(sig_B[20]), .B0(
        \mul/mult_6/n54 ), .B1(sig_B[19]), .C0(\mul/mult_6/n60 ), .C1(
        sig_B[18]), .Y(\mul/mult_6/n1082 ) );
  NAND2X2 \mul/mult_6/U1194  ( .A(sig_B[13]), .B(sig_B[14]), .Y(
        \mul/mult_6/n636 ) );
  NAND2X2 \mul/mult_6/U1147  ( .A(sig_B[18]), .B(sig_B[19]), .Y(
        \mul/mult_6/n604 ) );
  NAND2X2 \mul/mult_6/U1137  ( .A(sig_B[19]), .B(sig_B[20]), .Y(
        \mul/mult_6/n597 ) );
  NAND2X2 \mul/mult_6/U1129  ( .A(sig_B[20]), .B(sig_B[21]), .Y(
        \mul/mult_6/n592 ) );
  NAND2X2 \mul/mult_6/U1121  ( .A(sig_B[21]), .B(sig_B[22]), .Y(
        \mul/mult_6/n587 ) );
  AOI21X1 \mul/mult_6/U920  ( .A0(\mul/mult_6/n9 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n547 ), .Y(\mul/mult_6/n1338 ) );
  XOR2X1 \mul/mult_6/U464  ( .A(\mul/mult_6/n1014 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n774 ) );
  AOI21X1 \mul/mult_6/U837  ( .A0(\mul/mult_6/n20 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n543 ), .Y(\mul/mult_6/n1286 ) );
  AOI222XL \mul/mult_6/U537  ( .A0(n689), .A1(sig_B[14]), .B0(\mul/mult_6/n54 ), .B1(sig_B[13]), .C0(\mul/mult_6/n60 ), .C1(sig_B[12]), .Y(\mul/mult_6/n1088 ) );
  XOR2X1 \mul/mult_6/U461  ( .A(\mul/mult_6/n1013 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n773 ) );
  OAI21X1 \mul/mult_6/U459  ( .A0(n572), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1038 ), .Y(\mul/mult_6/n1012 ) );
  AOI222XL \mul/mult_6/U531  ( .A0(n689), .A1(sig_B[16]), .B0(\mul/mult_6/n54 ), .B1(sig_B[15]), .C0(\mul/mult_6/n60 ), .C1(sig_B[14]), .Y(\mul/mult_6/n1086 ) );
  AOI222XL \mul/mult_6/U682  ( .A0(\mul/mult_6/n32 ), .A1(sig_B[21]), .B0(n698), .B1(sig_B[20]), .C0(\mul/mult_6/n40 ), .C1(sig_B[19]), .Y(\mul/mult_6/n1185 ) );
  AOI222XL \mul/mult_6/U605  ( .A0(n687), .A1(sig_B[19]), .B0(n518), .B1(
        sig_B[18]), .C0(\mul/mult_6/n50 ), .C1(sig_B[17]), .Y(
        \mul/mult_6/n1135 ) );
  AOI222XL \mul/mult_6/U454  ( .A0(n692), .A1(sig_B[14]), .B0(\mul/mult_6/n64 ), .B1(sig_B[13]), .C0(\mul/mult_6/n70 ), .C1(sig_B[12]), .Y(\mul/mult_6/n1036 ) );
  AOI222XL \mul/mult_6/U528  ( .A0(n689), .A1(sig_B[17]), .B0(\mul/mult_6/n54 ), .B1(sig_B[16]), .C0(\mul/mult_6/n60 ), .C1(sig_B[15]), .Y(\mul/mult_6/n1085 ) );
  OAI21X1 \mul/mult_6/U674  ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1183 ), .Y(\mul/mult_6/n1157 ) );
  AOI222XL \mul/mult_6/U451  ( .A0(n692), .A1(sig_B[15]), .B0(\mul/mult_6/n64 ), .B1(sig_B[14]), .C0(\mul/mult_6/n70 ), .C1(sig_B[13]), .Y(\mul/mult_6/n1035 ) );
  OAI21X1 \mul/mult_6/U591  ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1131 ), .Y(\mul/mult_6/n1105 ) );
  NAND2XL \sigadd/add_9/U38  ( .A(n619), .B(\sigadd/add_9/n73 ), .Y(
        \sigadd/add_9/n6 ) );
  NAND2XL \sigadd/add_9/U52  ( .A(n593), .B(\sigadd/add_9/n81 ), .Y(
        \sigadd/add_9/n8 ) );
  NAND2BX2 \normal/srl_15/U246  ( .AN(n703), .B(add_out[48]), .Y(
        \normal/srl_15/n247 ) );
  AND3X6 \mul/mult_6/U1053  ( .A(\mul/mult_6/n1437 ), .B(\mul/mult_6/n1445 ), 
        .C(\mul/mult_6/n1453 ), .Y(\mul/mult_6/n70 ) );
  AO21X2 \mul/mult_6/U925  ( .A0(n701), .A1(sig_B[22]), .B0(n679), .Y(
        \mul/mult_6/n548 ) );
  AOI222XL \mul/mult_6/U703  ( .A0(n685), .A1(sig_B[14]), .B0(
        \mul/mult_6/n535 ), .B1(sig_B[13]), .C0(\mul/mult_6/n40 ), .C1(
        sig_B[12]), .Y(\mul/mult_6/n1192 ) );
  OAI21X1 \mul/mult_6/U702  ( .A0(n571), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1192 ), .Y(\mul/mult_6/n1166 ) );
  XOR2X1 \mul/mult_6/U479  ( .A(\mul/mult_6/n1019 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n779 ) );
  AOI222XL \mul/mult_6/U552  ( .A0(n689), .A1(sig_B[9]), .B0(n690), .B1(
        sig_B[8]), .C0(\mul/mult_6/n60 ), .C1(sig_B[7]), .Y(\mul/mult_6/n1093 ) );
  OAI21X1 \mul/mult_6/U551  ( .A0(n543), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1093 ), .Y(\mul/mult_6/n1067 ) );
  XOR2X1 \mul/mult_6/U550  ( .A(\mul/mult_6/n1067 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n802 ) );
  OAI21X1 \mul/mult_6/U625  ( .A0(n572), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1142 ), .Y(\mul/mult_6/n1116 ) );
  XOR2X1 \mul/mult_6/U624  ( .A(\mul/mult_6/n1116 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n826 ) );
  AOI222XL \mul/mult_6/U697  ( .A0(n685), .A1(sig_B[16]), .B0(
        \mul/mult_6/n535 ), .B1(sig_B[15]), .C0(\mul/mult_6/n40 ), .C1(
        sig_B[14]), .Y(\mul/mult_6/n1190 ) );
  OAI21X1 \mul/mult_6/U548  ( .A0(n542), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1092 ), .Y(\mul/mult_6/n1066 ) );
  XOR2X1 \mul/mult_6/U547  ( .A(\mul/mult_6/n1066 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n801 ) );
  XOR2X1 \mul/mult_6/U476  ( .A(\mul/mult_6/n1018 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n778 ) );
  XOR2X1 \mul/mult_6/U473  ( .A(\mul/mult_6/n1017 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n777 ) );
  AOI222XL \mul/mult_6/U700  ( .A0(n685), .A1(sig_B[15]), .B0(
        \mul/mult_6/n535 ), .B1(sig_B[14]), .C0(\mul/mult_6/n40 ), .C1(
        sig_B[13]), .Y(\mul/mult_6/n1191 ) );
  XOR2X1 \mul/mult_6/U627  ( .A(\mul/mult_6/n1117 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n827 ) );
  XOR2X1 \mul/mult_6/U918  ( .A(\mul/mult_6/n1312 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n922 ) );
  OAI21X1 \mul/mult_6/U622  ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1141 ), .Y(\mul/mult_6/n1115 ) );
  XOR2X1 \mul/mult_6/U621  ( .A(\mul/mult_6/n1115 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n825 ) );
  AOI21X1 \mul/mult_6/U841  ( .A0(\mul/mult_6/n20 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n544 ), .Y(\mul/mult_6/n1287 ) );
  XOR2X1 \mul/mult_6/U544  ( .A(\mul/mult_6/n1065 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n800 ) );
  OAI21X1 \mul/mult_6/U619  ( .A0(n571), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1140 ), .Y(\mul/mult_6/n1114 ) );
  XOR2X1 \mul/mult_6/U618  ( .A(\mul/mult_6/n1114 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n824 ) );
  XOR2X1 \mul/mult_6/U470  ( .A(\mul/mult_6/n1016 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n776 ) );
  AOI222XL \mul/mult_6/U768  ( .A0(\mul/mult_6/n22 ), .A1(sig_B[20]), .B0(n699), .B1(sig_B[19]), .C0(\mul/mult_6/n30 ), .C1(sig_B[18]), .Y(\mul/mult_6/n1238 ) );
  XOR2X1 \mul/mult_6/U766  ( .A(\mul/mult_6/n1212 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n872 ) );
  XOR2X1 \mul/mult_6/U832  ( .A(\mul/mult_6/n1259 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n894 ) );
  XOR2X1 \mul/mult_6/U541  ( .A(\mul/mult_6/n1064 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n799 ) );
  OAI21X1 \mul/mult_6/U468  ( .A0(n543), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1041 ), .Y(\mul/mult_6/n1015 ) );
  XOR2X1 \mul/mult_6/U467  ( .A(\mul/mult_6/n1015 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n775 ) );
  XOR2X1 \mul/mult_6/U689  ( .A(\mul/mult_6/n1162 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n847 ) );
  AOI222XL \mul/mult_6/U765  ( .A0(\mul/mult_6/n22 ), .A1(sig_B[21]), .B0(n699), .B1(sig_B[20]), .C0(\mul/mult_6/n30 ), .C1(sig_B[19]), .Y(\mul/mult_6/n1237 ) );
  XOR2X1 \mul/mult_6/U612  ( .A(\mul/mult_6/n1112 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n822 ) );
  AOI222XL \mul/mult_6/U617  ( .A0(n687), .A1(sig_B[15]), .B0(n518), .B1(
        sig_B[14]), .C0(\mul/mult_6/n50 ), .C1(sig_B[13]), .Y(
        \mul/mult_6/n1139 ) );
  XOR2X1 \mul/mult_6/U538  ( .A(\mul/mult_6/n1063 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n798 ) );
  AOI222XL \mul/mult_6/U762  ( .A0(\mul/mult_6/n22 ), .A1(sig_B[22]), .B0(n699), .B1(sig_B[21]), .C0(\mul/mult_6/n30 ), .C1(sig_B[20]), .Y(\mul/mult_6/n1236 ) );
  AOI21X1 \mul/mult_6/U758  ( .A0(\mul/mult_6/n30 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n540 ), .Y(\mul/mult_6/n1235 ) );
  AOI222XL \mul/mult_6/U460  ( .A0(n692), .A1(sig_B[12]), .B0(\mul/mult_6/n64 ), .B1(sig_B[11]), .C0(\mul/mult_6/n70 ), .C1(sig_B[10]), .Y(\mul/mult_6/n1038 ) );
  NAND2X2 \mul/mult_6/U1294  ( .A(sig_B[2]), .B(sig_B[3]), .Y(
        \mul/mult_6/n703 ) );
  NAND2X2 \mul/mult_6/U1269  ( .A(sig_B[5]), .B(sig_B[6]), .Y(
        \mul/mult_6/n687 ) );
  NOR2X2 \mul/mult_6/U1213  ( .A(sig_B[11]), .B(sig_B[12]), .Y(
        \mul/mult_6/n649 ) );
  NOR2X2 \mul/mult_6/U1193  ( .A(sig_B[13]), .B(sig_B[14]), .Y(
        \mul/mult_6/n635 ) );
  NAND2X2 \mul/mult_6/U1214  ( .A(sig_B[11]), .B(sig_B[12]), .Y(
        \mul/mult_6/n650 ) );
  NAND2X2 \mul/mult_6/U1186  ( .A(sig_B[14]), .B(sig_B[15]), .Y(
        \mul/mult_6/n631 ) );
  NAND2X2 \mul/mult_6/U1155  ( .A(sig_B[17]), .B(sig_B[18]), .Y(
        \mul/mult_6/n609 ) );
  AND3X6 \mul/mult_6/U1046  ( .A(\mul/mult_6/n1436 ), .B(\mul/mult_6/n1444 ), 
        .C(\mul/mult_6/n1452 ), .Y(\mul/mult_6/n78 ) );
  NAND2XL \sigadd/add_9/U66  ( .A(n594), .B(\sigadd/add_9/n89 ), .Y(
        \sigadd/add_9/n10 ) );
  NAND2X2 \mul/mult_6/U1233  ( .A(\mul/mult_6/n723 ), .B(\mul/mult_6/n666 ), 
        .Y(\mul/mult_6/n564 ) );
  ADDHX1 \mul/mult_6/U261  ( .A(\mul/mult_6/n386 ), .B(n609), .CO(
        \mul/mult_6/n375 ), .S(\mul/mult_6/n376 ) );
  AOI222XL \mul/mult_6/U789  ( .A0(n683), .A1(sig_B[13]), .B0(
        \mul/mult_6/n539 ), .B1(sig_B[12]), .C0(\mul/mult_6/n30 ), .C1(
        sig_B[11]), .Y(\mul/mult_6/n1245 ) );
  ADDHX1 \mul/mult_6/U257  ( .A(\mul/mult_6/n375 ), .B(n608), .CO(
        \mul/mult_6/n364 ), .S(\mul/mult_6/n365 ) );
  XOR2X1 \mul/mult_6/U559  ( .A(\mul/mult_6/n1070 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n805 ) );
  AOI222XL \mul/mult_6/U780  ( .A0(n683), .A1(sig_B[16]), .B0(
        \mul/mult_6/n539 ), .B1(sig_B[15]), .C0(\mul/mult_6/n30 ), .C1(
        sig_B[14]), .Y(\mul/mult_6/n1242 ) );
  XOR2X1 \mul/mult_6/U556  ( .A(\mul/mult_6/n1069 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n804 ) );
  AOI21X1 \mul/mult_6/U924  ( .A0(\mul/mult_6/n9 ), .A1(sig_B[21]), .B0(
        \mul/mult_6/n548 ), .Y(\mul/mult_6/n1339 ) );
  AOI222XL \mul/mult_6/U706  ( .A0(n685), .A1(sig_B[13]), .B0(
        \mul/mult_6/n535 ), .B1(sig_B[12]), .C0(\mul/mult_6/n40 ), .C1(
        sig_B[11]), .Y(\mul/mult_6/n1193 ) );
  OAI21X1 \mul/mult_6/U916  ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n8 ), 
        .B0(n680), .Y(\mul/mult_6/n1311 ) );
  OAI21X1 \mul/mult_6/U480  ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1045 ), .Y(\mul/mult_6/n1019 ) );
  AOI222XL \mul/mult_6/U774  ( .A0(n683), .A1(sig_B[18]), .B0(n699), .B1(
        sig_B[17]), .C0(\mul/mult_6/n30 ), .C1(sig_B[16]), .Y(
        \mul/mult_6/n1240 ) );
  XOR2X1 \mul/mult_6/U772  ( .A(\mul/mult_6/n1214 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n874 ) );
  AOI222XL \mul/mult_6/U848  ( .A0(\mul/mult_6/n12 ), .A1(sig_B[21]), .B0(n700), .B1(sig_B[20]), .C0(\mul/mult_6/n20 ), .C1(sig_B[19]), .Y(\mul/mult_6/n1289 ) );
  XOR2X1 \mul/mult_6/U846  ( .A(\mul/mult_6/n1263 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n898 ) );
  OAI21X1 \mul/mult_6/U477  ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1044 ), .Y(\mul/mult_6/n1018 ) );
  XOR2X1 \mul/mult_6/U698  ( .A(\mul/mult_6/n1165 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n850 ) );
  AOI222XL \mul/mult_6/U629  ( .A0(n687), .A1(sig_B[11]), .B0(n518), .B1(
        sig_B[10]), .C0(\mul/mult_6/n50 ), .C1(sig_B[9]), .Y(
        \mul/mult_6/n1143 ) );
  AOI222XL \mul/mult_6/U623  ( .A0(n687), .A1(sig_B[13]), .B0(n518), .B1(
        sig_B[12]), .C0(\mul/mult_6/n50 ), .C1(sig_B[11]), .Y(
        \mul/mult_6/n1141 ) );
  AOI222XL \mul/mult_6/U771  ( .A0(n683), .A1(sig_B[19]), .B0(n699), .B1(
        sig_B[18]), .C0(\mul/mult_6/n30 ), .C1(sig_B[17]), .Y(
        \mul/mult_6/n1239 ) );
  XOR2X1 \mul/mult_6/U769  ( .A(\mul/mult_6/n1213 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n873 ) );
  AOI222XL \mul/mult_6/U845  ( .A0(\mul/mult_6/n12 ), .A1(sig_B[22]), .B0(n700), .B1(sig_B[21]), .C0(\mul/mult_6/n20 ), .C1(sig_B[20]), .Y(\mul/mult_6/n1288 ) );
  XOR2X1 \mul/mult_6/U843  ( .A(\mul/mult_6/n1262 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n897 ) );
  XOR2X1 \mul/mult_6/U839  ( .A(\mul/mult_6/n1261 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n896 ) );
  AOI222XL \mul/mult_6/U694  ( .A0(n685), .A1(sig_B[17]), .B0(n698), .B1(
        sig_B[16]), .C0(\mul/mult_6/n40 ), .C1(sig_B[15]), .Y(
        \mul/mult_6/n1189 ) );
  XOR2X1 \mul/mult_6/U692  ( .A(\mul/mult_6/n1163 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n848 ) );
  AOI222XL \mul/mult_6/U620  ( .A0(n687), .A1(sig_B[14]), .B0(n518), .B1(
        sig_B[13]), .C0(\mul/mult_6/n50 ), .C1(sig_B[12]), .Y(
        \mul/mult_6/n1140 ) );
  OAI21X1 \mul/mult_6/U471  ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1042 ), .Y(\mul/mult_6/n1016 ) );
  OAI21X1 \mul/mult_6/U833  ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n18 ), 
        .B0(n682), .Y(\mul/mult_6/n1259 ) );
  AOI222XL \mul/mult_6/U469  ( .A0(n692), .A1(sig_B[9]), .B0(n693), .B1(
        sig_B[8]), .C0(\mul/mult_6/n70 ), .C1(sig_B[7]), .Y(\mul/mult_6/n1041 ) );
  XOR2X1 \mul/mult_6/U763  ( .A(\mul/mult_6/n1211 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n871 ) );
  XOR2X1 \mul/mult_6/U835  ( .A(\mul/mult_6/n1260 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n895 ) );
  OAI21X1 \mul/mult_6/U539  ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1089 ), .Y(\mul/mult_6/n1063 ) );
  AOI222XL \mul/mult_6/U688  ( .A0(n685), .A1(sig_B[19]), .B0(n698), .B1(
        sig_B[18]), .C0(\mul/mult_6/n40 ), .C1(sig_B[17]), .Y(
        \mul/mult_6/n1187 ) );
  XOR2X1 \mul/mult_6/U686  ( .A(\mul/mult_6/n1161 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n846 ) );
  XOR2X1 \mul/mult_6/U760  ( .A(\mul/mult_6/n1210 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n870 ) );
  XOR2X1 \mul/mult_6/U756  ( .A(\mul/mult_6/n1209 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n869 ) );
  XOR2X1 \mul/mult_6/U609  ( .A(\mul/mult_6/n1111 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n821 ) );
  OAI21X1 \mul/mult_6/U681  ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1185 ), .Y(\mul/mult_6/n1159 ) );
  OAI21X1 \mul/mult_6/U604  ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1135 ), .Y(\mul/mult_6/n1109 ) );
  OAI21X1 \mul/mult_6/U678  ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1184 ), .Y(\mul/mult_6/n1158 ) );
  OAI21X1 \mul/mult_6/U429  ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1028 ), .Y(\mul/mult_6/n1002 ) );
  NOR2X2 \mul/mult_6/U1284  ( .A(sig_B[3]), .B(sig_B[4]), .Y(\mul/mult_6/n696 ) );
  NAND2X2 \mul/mult_6/U1285  ( .A(sig_B[3]), .B(sig_B[4]), .Y(
        \mul/mult_6/n697 ) );
  NAND2X2 \mul/mult_6/U1263  ( .A(sig_B[6]), .B(sig_B[7]), .Y(
        \mul/mult_6/n684 ) );
  XNOR2X1 \mul/mult_6/U1092  ( .A(sig_A[3]), .B(sig_A[4]), .Y(
        \mul/mult_6/n1450 ) );
  NAND2XL \sigadd/add_9/U24  ( .A(n618), .B(\sigadd/add_9/n65 ), .Y(
        \sigadd/add_9/n4 ) );
  NAND2XL \sigadd/add_9/U58  ( .A(\sigadd/add_9/n255 ), .B(\sigadd/add_9/n84 ), 
        .Y(\sigadd/add_9/n9 ) );
  NAND2XL \sigadd/add_9/U72  ( .A(\sigadd/add_9/n257 ), .B(\sigadd/add_9/n92 ), 
        .Y(\sigadd/add_9/n11 ) );
  NAND2XL \sigadd/add_9/U80  ( .A(n595), .B(\sigadd/add_9/n97 ), .Y(
        \sigadd/add_9/n12 ) );
  NAND2XL \sigadd/add_9/U94  ( .A(n596), .B(\sigadd/add_9/n105 ), .Y(
        \sigadd/add_9/n14 ) );
  NAND2XL \sigadd/add_9/U108  ( .A(n597), .B(\sigadd/add_9/n113 ), .Y(
        \sigadd/add_9/n16 ) );
  NAND2X4 \round/r298/U116  ( .A(norm_out[9]), .B(norm_out[8]), .Y(
        \round/r298/n95 ) );
  NOR2X4 \ctrl/sub_0_root_add_0_root_sub_16/U45  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[1] ), .B(n710), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n33 ) );
  NAND2X2 \mul/mult_6/U1243  ( .A(\mul/mult_6/n724 ), .B(\mul/mult_6/n673 ), 
        .Y(\mul/mult_6/n565 ) );
  XNOR2X1 \mul/mult_6/U1071  ( .A(sig_A[12]), .B(sig_A[13]), .Y(
        \mul/mult_6/n1447 ) );
  ADDHX1 \mul/mult_6/U286  ( .A(sig_A[17]), .B(\mul/mult_6/n811 ), .CO(
        \mul/mult_6/n440 ), .S(\mul/mult_6/n441 ) );
  ADDHX1 \mul/mult_6/U273  ( .A(\mul/mult_6/n416 ), .B(\mul/mult_6/n783 ), 
        .CO(\mul/mult_6/n406 ), .S(\mul/mult_6/n407 ) );
  XOR2X1 \mul/mult_6/U784  ( .A(\mul/mult_6/n1218 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n878 ) );
  AOI222XL \mul/mult_6/U934  ( .A0(\mul/mult_6/n2 ), .A1(sig_B[20]), .B0(n701), 
        .B1(sig_B[19]), .C0(\mul/mult_6/n9 ), .C1(sig_B[18]), .Y(
        \mul/mult_6/n1342 ) );
  XOR2X1 \mul/mult_6/U932  ( .A(\mul/mult_6/n1316 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n926 ) );
  XOR2X1 \mul/mult_6/U787  ( .A(\mul/mult_6/n1219 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n879 ) );
  AOI222XL \mul/mult_6/U709  ( .A0(n685), .A1(sig_B[12]), .B0(
        \mul/mult_6/n535 ), .B1(sig_B[11]), .C0(\mul/mult_6/n40 ), .C1(
        sig_B[10]), .Y(\mul/mult_6/n1194 ) );
  XOR2X1 \mul/mult_6/U707  ( .A(\mul/mult_6/n1168 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n853 ) );
  OAI21X1 \mul/mult_6/U634  ( .A0(n543), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1145 ), .Y(\mul/mult_6/n1119 ) );
  AOI222XL \mul/mult_6/U783  ( .A0(n683), .A1(sig_B[15]), .B0(
        \mul/mult_6/n539 ), .B1(sig_B[14]), .C0(\mul/mult_6/n30 ), .C1(
        sig_B[13]), .Y(\mul/mult_6/n1243 ) );
  XOR2X1 \mul/mult_6/U781  ( .A(\mul/mult_6/n1217 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n877 ) );
  AOI222XL \mul/mult_6/U712  ( .A0(n685), .A1(sig_B[11]), .B0(
        \mul/mult_6/n535 ), .B1(sig_B[10]), .C0(\mul/mult_6/n40 ), .C1(
        sig_B[9]), .Y(\mul/mult_6/n1195 ) );
  XOR2X1 \mul/mult_6/U710  ( .A(\mul/mult_6/n1169 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n854 ) );
  AOI222XL \mul/mult_6/U931  ( .A0(\mul/mult_6/n2 ), .A1(sig_B[21]), .B0(n701), 
        .B1(sig_B[20]), .C0(\mul/mult_6/n9 ), .C1(sig_B[19]), .Y(
        \mul/mult_6/n1341 ) );
  XOR2X1 \mul/mult_6/U929  ( .A(\mul/mult_6/n1315 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n925 ) );
  OAI21X1 \mul/mult_6/U631  ( .A0(n542), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1144 ), .Y(\mul/mult_6/n1118 ) );
  OAI21X1 \mul/mult_6/U554  ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1094 ), .Y(\mul/mult_6/n1068 ) );
  XOR2X1 \mul/mult_6/U553  ( .A(\mul/mult_6/n1068 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n803 ) );
  AOI222XL \mul/mult_6/U777  ( .A0(n683), .A1(sig_B[17]), .B0(n699), .B1(
        sig_B[16]), .C0(\mul/mult_6/n30 ), .C1(sig_B[15]), .Y(
        \mul/mult_6/n1241 ) );
  XOR2X1 \mul/mult_6/U704  ( .A(\mul/mult_6/n1167 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n852 ) );
  AOI222XL \mul/mult_6/U928  ( .A0(\mul/mult_6/n2 ), .A1(sig_B[22]), .B0(n701), 
        .B1(sig_B[21]), .C0(\mul/mult_6/n9 ), .C1(sig_B[20]), .Y(
        \mul/mult_6/n1340 ) );
  OAI21X1 \mul/mult_6/U696  ( .A0(n570), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1190 ), .Y(\mul/mult_6/n1164 ) );
  OAI21X1 \mul/mult_6/U836  ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1286 ), .Y(\mul/mult_6/n1260 ) );
  NOR2X2 \mul/mult_6/U1227  ( .A(sig_B[10]), .B(sig_B[11]), .Y(
        \mul/mult_6/n660 ) );
  NAND2X2 \mul/mult_6/U1252  ( .A(sig_B[7]), .B(sig_B[8]), .Y(
        \mul/mult_6/n676 ) );
  NAND2X2 \mul/mult_6/U1173  ( .A(sig_B[15]), .B(sig_B[16]), .Y(
        \mul/mult_6/n621 ) );
  AOI222XL \mul/mult_6/U896  ( .A0(n681), .A1(sig_B[5]), .B0(\mul/mult_6/n543 ), .B1(sig_B[4]), .C0(\mul/mult_6/n20 ), .C1(sig_B[3]), .Y(\mul/mult_6/n1305 )
         );
  NAND2X2 \sigadd/add_9/U41  ( .A(ali_P[44]), .B(ali_C[44]), .Y(
        \sigadd/add_9/n73 ) );
  NAND2XL \sigadd/add_9/U86  ( .A(\sigadd/add_9/n259 ), .B(\sigadd/add_9/n100 ), .Y(\sigadd/add_9/n13 ) );
  NAND2XL \sigadd/add_9/U100  ( .A(\sigadd/add_9/n261 ), .B(
        \sigadd/add_9/n108 ), .Y(\sigadd/add_9/n15 ) );
  NAND2XL \sigadd/add_9/U122  ( .A(n598), .B(\sigadd/add_9/n121 ), .Y(
        \sigadd/add_9/n18 ) );
  NAND2XL \sigadd/add_9/U136  ( .A(n599), .B(\sigadd/add_9/n129 ), .Y(
        \sigadd/add_9/n20 ) );
  NAND2XL \sigadd/add_9/U150  ( .A(n573), .B(\sigadd/add_9/n137 ), .Y(
        \sigadd/add_9/n22 ) );
  XNOR2X1 \mul/mult_6/U1078  ( .A(sig_A[9]), .B(sig_A[10]), .Y(
        \mul/mult_6/n1448 ) );
  AND3X6 \mul/mult_6/U1060  ( .A(\mul/mult_6/n1438 ), .B(\mul/mult_6/n1446 ), 
        .C(\mul/mult_6/n1454 ), .Y(\mul/mult_6/n60 ) );
  ADDHX1 \mul/mult_6/U283  ( .A(\mul/mult_6/n440 ), .B(\mul/mult_6/n810 ), 
        .CO(\mul/mult_6/n432 ), .S(\mul/mult_6/n433 ) );
  XOR2X1 \mul/mult_6/U565  ( .A(\mul/mult_6/n1072 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n807 ) );
  AOI222XL \mul/mult_6/U875  ( .A0(n681), .A1(sig_B[12]), .B0(
        \mul/mult_6/n543 ), .B1(sig_B[11]), .C0(\mul/mult_6/n20 ), .C1(
        sig_B[10]), .Y(\mul/mult_6/n1298 ) );
  AOI222XL \mul/mult_6/U801  ( .A0(n683), .A1(sig_B[9]), .B0(\mul/mult_6/n539 ), .B1(sig_B[8]), .C0(\mul/mult_6/n30 ), .C1(sig_B[7]), .Y(\mul/mult_6/n1249 )
         );
  AOI222XL \mul/mult_6/U798  ( .A0(n683), .A1(sig_B[10]), .B0(
        \mul/mult_6/n539 ), .B1(sig_B[9]), .C0(\mul/mult_6/n30 ), .C1(sig_B[8]), .Y(\mul/mult_6/n1248 ) );
  AOI222XL \mul/mult_6/U724  ( .A0(n685), .A1(sig_B[7]), .B0(\mul/mult_6/n535 ), .B1(sig_B[6]), .C0(\mul/mult_6/n40 ), .C1(sig_B[5]), .Y(\mul/mult_6/n1199 )
         );
  XOR2X1 \mul/mult_6/U719  ( .A(\mul/mult_6/n1172 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n857 ) );
  AOI222XL \mul/mult_6/U869  ( .A0(n681), .A1(sig_B[14]), .B0(
        \mul/mult_6/n543 ), .B1(sig_B[13]), .C0(\mul/mult_6/n20 ), .C1(
        sig_B[12]), .Y(\mul/mult_6/n1296 ) );
  AOI222XL \mul/mult_6/U792  ( .A0(n683), .A1(sig_B[12]), .B0(
        \mul/mult_6/n539 ), .B1(sig_B[11]), .C0(\mul/mult_6/n30 ), .C1(
        sig_B[10]), .Y(\mul/mult_6/n1246 ) );
  AOI222XL \mul/mult_6/U795  ( .A0(n683), .A1(sig_B[11]), .B0(
        \mul/mult_6/n539 ), .B1(sig_B[10]), .C0(\mul/mult_6/n30 ), .C1(
        sig_B[9]), .Y(\mul/mult_6/n1247 ) );
  XOR2X1 \mul/mult_6/U793  ( .A(\mul/mult_6/n1221 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n881 ) );
  AOI222XL \mul/mult_6/U863  ( .A0(n681), .A1(sig_B[16]), .B0(
        \mul/mult_6/n543 ), .B1(sig_B[15]), .C0(\mul/mult_6/n20 ), .C1(
        sig_B[14]), .Y(\mul/mult_6/n1294 ) );
  XOR2X1 \mul/mult_6/U636  ( .A(\mul/mult_6/n1120 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n830 ) );
  XOR2X1 \mul/mult_6/U562  ( .A(\mul/mult_6/n1071 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n806 ) );
  AOI222XL \mul/mult_6/U866  ( .A0(n681), .A1(sig_B[15]), .B0(
        \mul/mult_6/n543 ), .B1(sig_B[14]), .C0(\mul/mult_6/n20 ), .C1(
        sig_B[13]), .Y(\mul/mult_6/n1295 ) );
  XOR2X1 \mul/mult_6/U935  ( .A(\mul/mult_6/n1317 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n927 ) );
  XOR2X1 \mul/mult_6/U855  ( .A(\mul/mult_6/n1266 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n901 ) );
  AOI222XL \mul/mult_6/U860  ( .A0(\mul/mult_6/n12 ), .A1(sig_B[17]), .B0(n700), .B1(sig_B[16]), .C0(\mul/mult_6/n20 ), .C1(sig_B[15]), .Y(\mul/mult_6/n1293 ) );
  XOR2X1 \mul/mult_6/U858  ( .A(\mul/mult_6/n1267 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n902 ) );
  AOI222XL \mul/mult_6/U635  ( .A0(n687), .A1(sig_B[9]), .B0(n518), .B1(
        sig_B[8]), .C0(\mul/mult_6/n50 ), .C1(sig_B[7]), .Y(\mul/mult_6/n1145 ) );
  AOI222XL \mul/mult_6/U632  ( .A0(n687), .A1(sig_B[10]), .B0(n518), .B1(
        sig_B[9]), .C0(\mul/mult_6/n50 ), .C1(sig_B[8]), .Y(\mul/mult_6/n1144 ) );
  XOR2X1 \mul/mult_6/U778  ( .A(\mul/mult_6/n1216 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n876 ) );
  AOI222XL \mul/mult_6/U851  ( .A0(\mul/mult_6/n12 ), .A1(sig_B[20]), .B0(n700), .B1(sig_B[19]), .C0(\mul/mult_6/n20 ), .C1(sig_B[18]), .Y(\mul/mult_6/n1290 ) );
  XOR2X1 \mul/mult_6/U849  ( .A(\mul/mult_6/n1264 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n899 ) );
  XOR2X1 \mul/mult_6/U922  ( .A(\mul/mult_6/n1313 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n923 ) );
  XOR2X1 \mul/mult_6/U775  ( .A(\mul/mult_6/n1215 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n875 ) );
  XOR2X1 \mul/mult_6/U926  ( .A(\mul/mult_6/n1314 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n924 ) );
  OAI21X1 \mul/mult_6/U773  ( .A0(n569), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1240 ), .Y(\mul/mult_6/n1214 ) );
  AOI222XL \mul/mult_6/U475  ( .A0(n692), .A1(sig_B[7]), .B0(n693), .B1(
        sig_B[6]), .C0(\mul/mult_6/n70 ), .C1(sig_B[5]), .Y(\mul/mult_6/n1043 ) );
  OAI21X1 \mul/mult_6/U699  ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1191 ), .Y(\mul/mult_6/n1165 ) );
  OAI21X1 \mul/mult_6/U628  ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1143 ), .Y(\mul/mult_6/n1117 ) );
  OAI21X1 \mul/mult_6/U767  ( .A0(n591), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1238 ), .Y(\mul/mult_6/n1212 ) );
  OAI21X1 \mul/mult_6/U690  ( .A0(n569), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1188 ), .Y(\mul/mult_6/n1162 ) );
  OAI21X1 \mul/mult_6/U616  ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1139 ), .Y(\mul/mult_6/n1113 ) );
  AOI222XL \mul/mult_6/U540  ( .A0(n689), .A1(sig_B[13]), .B0(n690), .B1(
        sig_B[12]), .C0(\mul/mult_6/n60 ), .C1(sig_B[11]), .Y(
        \mul/mult_6/n1089 ) );
  NOR2X2 \mul/mult_6/U1289  ( .A(\mul/mult_6/n705 ), .B(\mul/mult_6/n702 ), 
        .Y(\mul/mult_6/n700 ) );
  NOR2X2 \mul/mult_6/U1272  ( .A(\mul/mult_6/n696 ), .B(\mul/mult_6/n691 ), 
        .Y(\mul/mult_6/n689 ) );
  NAND2X2 \mul/mult_6/U1246  ( .A(sig_B[8]), .B(sig_B[9]), .Y(
        \mul/mult_6/n673 ) );
  OAI21X1 \mul/mult_6/U1143  ( .A0(\mul/mult_6/n603 ), .A1(\mul/mult_6/n609 ), 
        .B0(\mul/mult_6/n604 ), .Y(\mul/mult_6/n602 ) );
  MXI2X2 \align/sra_10/U258  ( .A(\align/sra_10/n296 ), .B(\align/sra_10/n297 ), .S0(n507), .Y(\align/sra_10/n242 ) );
  NAND2X2 \sigadd/add_9/U27  ( .A(ali_P[46]), .B(ali_C[46]), .Y(
        \sigadd/add_9/n65 ) );
  NAND2X2 \sigadd/add_9/U13  ( .A(ali_P[48]), .B(ali_C[48]), .Y(
        \sigadd/add_9/n57 ) );
  NAND2XL \sigadd/add_9/U44  ( .A(\sigadd/add_9/n253 ), .B(\sigadd/add_9/n76 ), 
        .Y(\sigadd/add_9/n7 ) );
  NAND2XL \sigadd/add_9/U114  ( .A(\sigadd/add_9/n263 ), .B(
        \sigadd/add_9/n116 ), .Y(\sigadd/add_9/n17 ) );
  NAND2XL \sigadd/add_9/U128  ( .A(\sigadd/add_9/n265 ), .B(
        \sigadd/add_9/n124 ), .Y(\sigadd/add_9/n19 ) );
  NAND2XL \sigadd/add_9/U164  ( .A(n574), .B(\sigadd/add_9/n145 ), .Y(
        \sigadd/add_9/n24 ) );
  NAND2XL \sigadd/add_9/U178  ( .A(n575), .B(\sigadd/add_9/n153 ), .Y(
        \sigadd/add_9/n26 ) );
  NAND2XL \sigadd/add_9/U10  ( .A(n617), .B(\sigadd/add_9/n57 ), .Y(
        \sigadd/add_9/n2 ) );
  ADDHX1 \mul/mult_6/U292  ( .A(\mul/mult_6/n461 ), .B(\mul/mult_6/n837 ), 
        .CO(\mul/mult_6/n454 ), .S(\mul/mult_6/n455 ) );
  XOR2X1 \mul/mult_6/U578  ( .A(\mul/mult_6/n1076 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n811 ) );
  AOI222XL \mul/mult_6/U807  ( .A0(n683), .A1(sig_B[7]), .B0(\mul/mult_6/n539 ), .B1(sig_B[6]), .C0(\mul/mult_6/n30 ), .C1(sig_B[5]), .Y(\mul/mult_6/n1251 )
         );
  NAND2X2 \mul/mult_6/U1197  ( .A(\mul/mult_6/n654 ), .B(\mul/mult_6/n640 ), 
        .Y(\mul/mult_6/n638 ) );
  AOI222XL \mul/mult_6/U727  ( .A0(n685), .A1(sig_B[6]), .B0(\mul/mult_6/n535 ), .B1(sig_B[5]), .C0(\mul/mult_6/n40 ), .C1(sig_B[4]), .Y(\mul/mult_6/n1200 )
         );
  OAI21X1 \mul/mult_6/U649  ( .A0(n545), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1150 ), .Y(\mul/mult_6/n1124 ) );
  XOR2X1 \mul/mult_6/U799  ( .A(\mul/mult_6/n1223 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n883 ) );
  AOI222XL \mul/mult_6/U946  ( .A0(n679), .A1(sig_B[16]), .B0(
        \mul/mult_6/n547 ), .B1(sig_B[15]), .C0(\mul/mult_6/n9 ), .C1(
        sig_B[14]), .Y(\mul/mult_6/n1346 ) );
  OAI21X1 \mul/mult_6/U646  ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1149 ), .Y(\mul/mult_6/n1123 ) );
  AOI222XL \mul/mult_6/U721  ( .A0(n685), .A1(sig_B[8]), .B0(\mul/mult_6/n535 ), .B1(sig_B[7]), .C0(\mul/mult_6/n40 ), .C1(sig_B[6]), .Y(\mul/mult_6/n1198 )
         );
  OAI21X1 \mul/mult_6/U720  ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1198 ), .Y(\mul/mult_6/n1172 ) );
  AOI222XL \mul/mult_6/U872  ( .A0(n681), .A1(sig_B[13]), .B0(
        \mul/mult_6/n543 ), .B1(sig_B[12]), .C0(\mul/mult_6/n20 ), .C1(
        sig_B[11]), .Y(\mul/mult_6/n1297 ) );
  XOR2X1 \mul/mult_6/U870  ( .A(\mul/mult_6/n1271 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n906 ) );
  AOI222XL \mul/mult_6/U718  ( .A0(n685), .A1(sig_B[9]), .B0(\mul/mult_6/n535 ), .B1(sig_B[8]), .C0(\mul/mult_6/n40 ), .C1(sig_B[7]), .Y(\mul/mult_6/n1197 )
         );
  OAI21X1 \mul/mult_6/U717  ( .A0(n543), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1197 ), .Y(\mul/mult_6/n1171 ) );
  XOR2X1 \mul/mult_6/U716  ( .A(\mul/mult_6/n1171 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n856 ) );
  AOI222XL \mul/mult_6/U715  ( .A0(n685), .A1(sig_B[10]), .B0(
        \mul/mult_6/n535 ), .B1(sig_B[9]), .C0(\mul/mult_6/n40 ), .C1(sig_B[8]), .Y(\mul/mult_6/n1196 ) );
  XOR2X1 \mul/mult_6/U713  ( .A(\mul/mult_6/n1170 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n855 ) );
  OAI21X1 \mul/mult_6/U640  ( .A0(n544), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1147 ), .Y(\mul/mult_6/n1121 ) );
  OAI21X1 \mul/mult_6/U785  ( .A0(n571), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1244 ), .Y(\mul/mult_6/n1218 ) );
  AOI222XL \mul/mult_6/U937  ( .A0(n679), .A1(sig_B[19]), .B0(n701), .B1(
        sig_B[18]), .C0(\mul/mult_6/n9 ), .C1(sig_B[17]), .Y(
        \mul/mult_6/n1343 ) );
  OAI21X1 \mul/mult_6/U788  ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1245 ), .Y(\mul/mult_6/n1219 ) );
  AOI222XL \mul/mult_6/U407  ( .A0(n695), .A1(sig_B[2]), .B0(n696), .B1(
        sig_B[1]), .C0(\mul/mult_6/n78 ), .C1(sig_B[0]), .Y(\mul/mult_6/n996 )
         );
  OAI21X1 \mul/mult_6/U708  ( .A0(n572), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1194 ), .Y(\mul/mult_6/n1168 ) );
  AOI222XL \mul/mult_6/U857  ( .A0(n681), .A1(sig_B[18]), .B0(n700), .B1(
        sig_B[17]), .C0(\mul/mult_6/n20 ), .C1(sig_B[16]), .Y(
        \mul/mult_6/n1292 ) );
  OAI21X1 \mul/mult_6/U711  ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1195 ), .Y(\mul/mult_6/n1169 ) );
  OAI21X1 \mul/mult_6/U705  ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1193 ), .Y(\mul/mult_6/n1167 ) );
  XOR2X1 \mul/mult_6/U852  ( .A(\mul/mult_6/n1265 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n900 ) );
  AOI222XL \mul/mult_6/U481  ( .A0(n692), .A1(sig_B[5]), .B0(\mul/mult_6/n64 ), 
        .B1(sig_B[4]), .C0(\mul/mult_6/n70 ), .C1(sig_B[3]), .Y(
        \mul/mult_6/n1045 ) );
  AOI222XL \mul/mult_6/U549  ( .A0(n689), .A1(sig_B[10]), .B0(n690), .B1(
        sig_B[9]), .C0(\mul/mult_6/n60 ), .C1(sig_B[8]), .Y(\mul/mult_6/n1092 ) );
  AOI222XL \mul/mult_6/U478  ( .A0(n692), .A1(sig_B[6]), .B0(n693), .B1(
        sig_B[5]), .C0(\mul/mult_6/n70 ), .C1(sig_B[4]), .Y(\mul/mult_6/n1044 ) );
  AOI222XL \mul/mult_6/U398  ( .A0(n695), .A1(sig_B[5]), .B0(n696), .B1(
        sig_B[4]), .C0(\mul/mult_6/n78 ), .C1(sig_B[3]), .Y(\mul/mult_6/n993 )
         );
  OAI21X1 \mul/mult_6/U770  ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1239 ), .Y(\mul/mult_6/n1213 ) );
  OAI21X1 \mul/mult_6/U693  ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1189 ), .Y(\mul/mult_6/n1163 ) );
  AOI222XL \mul/mult_6/U395  ( .A0(n695), .A1(sig_B[6]), .B0(n696), .B1(
        sig_B[5]), .C0(\mul/mult_6/n78 ), .C1(sig_B[4]), .Y(\mul/mult_6/n992 )
         );
  OAI21X1 \mul/mult_6/U764  ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1237 ), .Y(\mul/mult_6/n1211 ) );
  OAI21X1 \mul/mult_6/U687  ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1187 ), .Y(\mul/mult_6/n1161 ) );
  AND3X6 \mul/mult_6/U1081  ( .A(\mul/mult_6/n1441 ), .B(\mul/mult_6/n1449 ), 
        .C(\mul/mult_6/n1457 ), .Y(\mul/mult_6/n30 ) );
  OAI21X1 \mul/mult_6/U969  ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1354 ), .Y(\mul/mult_6/n1328 ) );
  AOI222XL \mul/mult_6/U973  ( .A0(n679), .A1(sig_B[7]), .B0(\mul/mult_6/n547 ), .B1(sig_B[6]), .C0(\mul/mult_6/n9 ), .C1(sig_B[5]), .Y(\mul/mult_6/n1355 )
         );
  MXI2X2 \align/sra_10/U262  ( .A(\align/sra_10/n292 ), .B(\align/sra_10/n293 ), .S0(n507), .Y(\align/sra_10/n238 ) );
  MXI2X2 \align/sra_10/U260  ( .A(\align/sra_10/n294 ), .B(\align/sra_10/n295 ), .S0(n507), .Y(\align/sra_10/n240 ) );
  NAND2XL \sigadd/add_9/U142  ( .A(\sigadd/add_9/n267 ), .B(
        \sigadd/add_9/n132 ), .Y(\sigadd/add_9/n21 ) );
  NAND2XL \sigadd/add_9/U156  ( .A(\sigadd/add_9/n269 ), .B(
        \sigadd/add_9/n140 ), .Y(\sigadd/add_9/n23 ) );
  NAND2XL \sigadd/add_9/U170  ( .A(\sigadd/add_9/n271 ), .B(
        \sigadd/add_9/n148 ), .Y(\sigadd/add_9/n25 ) );
  NAND2XL \sigadd/add_9/U184  ( .A(\sigadd/add_9/n273 ), .B(
        \sigadd/add_9/n156 ), .Y(\sigadd/add_9/n27 ) );
  NAND2XL \sigadd/add_9/U192  ( .A(n576), .B(\sigadd/add_9/n161 ), .Y(
        \sigadd/add_9/n28 ) );
  NAND2XL \sigadd/add_9/U206  ( .A(n577), .B(\sigadd/add_9/n169 ), .Y(
        \sigadd/add_9/n30 ) );
  NAND2XL \sigadd/add_9/U220  ( .A(n578), .B(\sigadd/add_9/n177 ), .Y(
        \sigadd/add_9/n32 ) );
  NAND2XL \sigadd/add_9/U16  ( .A(\sigadd/add_9/n249 ), .B(\sigadd/add_9/n60 ), 
        .Y(\sigadd/add_9/n3 ) );
  AND3X6 \mul/mult_6/U1074  ( .A(\mul/mult_6/n1440 ), .B(\mul/mult_6/n1448 ), 
        .C(\mul/mult_6/n1456 ), .Y(\mul/mult_6/n40 ) );
  AOI222XL \mul/mult_6/U804  ( .A0(n683), .A1(sig_B[8]), .B0(\mul/mult_6/n539 ), .B1(sig_B[7]), .C0(\mul/mult_6/n30 ), .C1(sig_B[6]), .Y(\mul/mult_6/n1250 )
         );
  AOI222XL \mul/mult_6/U730  ( .A0(n685), .A1(sig_B[5]), .B0(\mul/mult_6/n535 ), .B1(sig_B[4]), .C0(\mul/mult_6/n40 ), .C1(sig_B[3]), .Y(\mul/mult_6/n1201 )
         );
  AOI222XL \mul/mult_6/U813  ( .A0(n683), .A1(sig_B[5]), .B0(\mul/mult_6/n539 ), .B1(sig_B[4]), .C0(\mul/mult_6/n30 ), .C1(sig_B[3]), .Y(\mul/mult_6/n1253 )
         );
  AOI222XL \mul/mult_6/U810  ( .A0(n683), .A1(sig_B[6]), .B0(\mul/mult_6/n539 ), .B1(sig_B[5]), .C0(\mul/mult_6/n30 ), .C1(sig_B[4]), .Y(\mul/mult_6/n1252 )
         );
  AOI222XL \mul/mult_6/U884  ( .A0(n681), .A1(sig_B[9]), .B0(\mul/mult_6/n543 ), .B1(sig_B[8]), .C0(\mul/mult_6/n20 ), .C1(sig_B[7]), .Y(\mul/mult_6/n1301 )
         );
  AOI222XL \mul/mult_6/U881  ( .A0(n681), .A1(sig_B[10]), .B0(
        \mul/mult_6/n543 ), .B1(sig_B[9]), .C0(\mul/mult_6/n20 ), .C1(sig_B[8]), .Y(\mul/mult_6/n1300 ) );
  XOR2X1 \mul/mult_6/U879  ( .A(\mul/mult_6/n1274 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n909 ) );
  XOR2X1 \mul/mult_6/U574  ( .A(\mul/mult_6/n1075 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n810 ) );
  XOR2X1 \mul/mult_6/U568  ( .A(\mul/mult_6/n1073 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n808 ) );
  ADDFX1 \mul/mult_6/U276  ( .A(\mul/mult_6/n417 ), .B(\mul/mult_6/n808 ), 
        .CI(\mul/mult_6/n424 ), .CO(\mul/mult_6/n414 ), .S(\mul/mult_6/n415 )
         );
  AOI222XL \mul/mult_6/U878  ( .A0(n681), .A1(sig_B[11]), .B0(
        \mul/mult_6/n543 ), .B1(sig_B[10]), .C0(\mul/mult_6/n20 ), .C1(
        sig_B[9]), .Y(\mul/mult_6/n1299 ) );
  OAI21X1 \mul/mult_6/U800  ( .A0(n543), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1249 ), .Y(\mul/mult_6/n1223 ) );
  AOI222XL \mul/mult_6/U949  ( .A0(n679), .A1(sig_B[15]), .B0(
        \mul/mult_6/n547 ), .B1(sig_B[14]), .C0(\mul/mult_6/n9 ), .C1(
        sig_B[13]), .Y(\mul/mult_6/n1347 ) );
  OAI21X1 \mul/mult_6/U723  ( .A0(n544), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1199 ), .Y(\mul/mult_6/n1173 ) );
  AOI222XL \mul/mult_6/U943  ( .A0(n679), .A1(sig_B[17]), .B0(n701), .B1(
        sig_B[16]), .C0(\mul/mult_6/n9 ), .C1(sig_B[15]), .Y(
        \mul/mult_6/n1345 ) );
  XOR2X1 \mul/mult_6/U941  ( .A(\mul/mult_6/n1319 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n929 ) );
  XOR2X1 \mul/mult_6/U861  ( .A(\mul/mult_6/n1268 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n903 ) );
  OAI21X1 \mul/mult_6/U637  ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1146 ), .Y(\mul/mult_6/n1120 ) );
  AOI222XL \mul/mult_6/U940  ( .A0(n679), .A1(sig_B[18]), .B0(n701), .B1(
        sig_B[17]), .C0(\mul/mult_6/n9 ), .C1(sig_B[16]), .Y(
        \mul/mult_6/n1344 ) );
  XOR2X1 \mul/mult_6/U938  ( .A(\mul/mult_6/n1318 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n928 ) );
  XOR2X1 \mul/mult_6/U864  ( .A(\mul/mult_6/n1269 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n904 ) );
  OAI21X1 \mul/mult_6/U779  ( .A0(n570), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1242 ), .Y(\mul/mult_6/n1216 ) );
  AOI222XL \mul/mult_6/U558  ( .A0(n689), .A1(sig_B[7]), .B0(n690), .B1(
        sig_B[6]), .C0(\mul/mult_6/n60 ), .C1(sig_B[5]), .Y(\mul/mult_6/n1095 ) );
  OAI21X1 \mul/mult_6/U850  ( .A0(n591), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1290 ), .Y(\mul/mult_6/n1264 ) );
  AOI222XL \mul/mult_6/U854  ( .A0(\mul/mult_6/n12 ), .A1(sig_B[19]), .B0(n700), .B1(sig_B[18]), .C0(\mul/mult_6/n20 ), .C1(sig_B[17]), .Y(\mul/mult_6/n1291 ) );
  AOI222XL \mul/mult_6/U626  ( .A0(n687), .A1(sig_B[12]), .B0(n518), .B1(
        sig_B[11]), .C0(\mul/mult_6/n50 ), .C1(sig_B[10]), .Y(
        \mul/mult_6/n1142 ) );
  OAI21X1 \mul/mult_6/U847  ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1289 ), .Y(\mul/mult_6/n1263 ) );
  OAI21X1 \mul/mult_6/U844  ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1288 ), .Y(\mul/mult_6/n1262 ) );
  OAI21X1 \mul/mult_6/U761  ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1236 ), .Y(\mul/mult_6/n1210 ) );
  ADDFX1 \expadd/add_0_root_sub_0_root_sub_8/U7  ( .A(\expadd/N2 ), .B(
        exp_B[2]), .CI(\expadd/add_0_root_sub_0_root_sub_8/n8 ), .CO(
        \expadd/add_0_root_sub_0_root_sub_8/n7 ), .S(exp_P[2]) );
  ADDFX1 \expadd/add_0_root_sub_0_root_sub_8/U8  ( .A(
        \expadd/add_0_root_sub_0_root_sub_8/n9 ), .B(exp_B[1]), .CI(
        \expadd/N1 ), .CO(\expadd/add_0_root_sub_0_root_sub_8/n8 ), .S(
        exp_P[1]) );
  NAND2X2 \mul/mult_6/U1300  ( .A(sig_B[1]), .B(sig_B[2]), .Y(
        \mul/mult_6/n706 ) );
  NOR2X2 \mul/mult_6/U1268  ( .A(sig_B[5]), .B(sig_B[6]), .Y(\mul/mult_6/n686 ) );
  CLKXOR2X2 \mul/mult_6/U1087  ( .A(sig_A[7]), .B(sig_A[8]), .Y(
        \mul/mult_6/n1457 ) );
  XNOR2X1 \mul/mult_6/U1085  ( .A(sig_A[6]), .B(sig_A[7]), .Y(
        \mul/mult_6/n1449 ) );
  XOR2X1 \mul/mult_6/U1247  ( .A(\mul/mult_6/n677 ), .B(\mul/mult_6/n566 ), 
        .Y(\mul/mult_6/n1405 ) );
  XOR2X1 \mul/mult_6/U1270  ( .A(\mul/mult_6/n693 ), .B(\mul/mult_6/n569 ), 
        .Y(\mul/mult_6/n1408 ) );
  MXI2X2 \align/sra_10/U266  ( .A(\align/sra_10/n288 ), .B(\align/sra_10/n289 ), .S0(n507), .Y(\align/sra_10/n234 ) );
  MXI2X2 \align/sra_10/U264  ( .A(\align/sra_10/n290 ), .B(\align/sra_10/n291 ), .S0(n507), .Y(\align/sra_10/n236 ) );
  NAND2XL \sigadd/add_9/U198  ( .A(\sigadd/add_9/n275 ), .B(
        \sigadd/add_9/n164 ), .Y(\sigadd/add_9/n29 ) );
  NAND2XL \sigadd/add_9/U212  ( .A(\sigadd/add_9/n277 ), .B(
        \sigadd/add_9/n172 ), .Y(\sigadd/add_9/n31 ) );
  NAND2XL \sigadd/add_9/U226  ( .A(\sigadd/add_9/n279 ), .B(
        \sigadd/add_9/n180 ), .Y(\sigadd/add_9/n33 ) );
  NAND2XL \sigadd/add_9/U234  ( .A(n579), .B(\sigadd/add_9/n185 ), .Y(
        \sigadd/add_9/n34 ) );
  NAND2XL \sigadd/add_9/U248  ( .A(n547), .B(\sigadd/add_9/n193 ), .Y(
        \sigadd/add_9/n36 ) );
  OAI21X1 \mul/mult_6/U732  ( .A0(n545), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1202 ), .Y(\mul/mult_6/n1176 ) );
  ADDFX1 \mul/mult_6/U294  ( .A(\mul/mult_6/n462 ), .B(\mul/mult_6/n862 ), 
        .CI(\mul/mult_6/n466 ), .CO(\mul/mult_6/n459 ), .S(\mul/mult_6/n460 )
         );
  ADDFX1 \mul/mult_6/U291  ( .A(\mul/mult_6/n455 ), .B(\mul/mult_6/n861 ), 
        .CI(\mul/mult_6/n459 ), .CO(\mul/mult_6/n452 ), .S(\mul/mult_6/n453 )
         );
  ADDHX1 \mul/mult_6/U289  ( .A(\mul/mult_6/n836 ), .B(\mul/mult_6/n454 ), 
        .CO(\mul/mult_6/n447 ), .S(\mul/mult_6/n448 ) );
  XOR2X1 \mul/mult_6/U885  ( .A(\mul/mult_6/n1276 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n911 ) );
  ADDFX1 \mul/mult_6/U288  ( .A(\mul/mult_6/n448 ), .B(\mul/mult_6/n884 ), 
        .CI(\mul/mult_6/n860 ), .CO(\mul/mult_6/n445 ), .S(\mul/mult_6/n446 )
         );
  AOI222XL \mul/mult_6/U958  ( .A0(n679), .A1(sig_B[12]), .B0(
        \mul/mult_6/n547 ), .B1(sig_B[11]), .C0(\mul/mult_6/n9 ), .C1(
        sig_B[10]), .Y(\mul/mult_6/n1350 ) );
  AOI222XL \mul/mult_6/U961  ( .A0(n679), .A1(sig_B[11]), .B0(
        \mul/mult_6/n547 ), .B1(sig_B[10]), .C0(\mul/mult_6/n9 ), .C1(sig_B[9]), .Y(\mul/mult_6/n1351 ) );
  XOR2X1 \mul/mult_6/U571  ( .A(\mul/mult_6/n1074 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n809 ) );
  AOI222XL \mul/mult_6/U955  ( .A0(n679), .A1(sig_B[13]), .B0(
        \mul/mult_6/n547 ), .B1(sig_B[12]), .C0(\mul/mult_6/n9 ), .C1(
        sig_B[11]), .Y(\mul/mult_6/n1349 ) );
  AOI222XL \mul/mult_6/U952  ( .A0(n679), .A1(sig_B[14]), .B0(
        \mul/mult_6/n547 ), .B1(sig_B[13]), .C0(\mul/mult_6/n9 ), .C1(
        sig_B[12]), .Y(\mul/mult_6/n1348 ) );
  OAI21X1 \mul/mult_6/U874  ( .A0(n572), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1298 ), .Y(\mul/mult_6/n1272 ) );
  OAI21X1 \mul/mult_6/U797  ( .A0(n542), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1248 ), .Y(\mul/mult_6/n1222 ) );
  OAI21X1 \mul/mult_6/U791  ( .A0(n572), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1246 ), .Y(\mul/mult_6/n1220 ) );
  OAI21X1 \mul/mult_6/U714  ( .A0(n542), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1196 ), .Y(\mul/mult_6/n1170 ) );
  AOI222XL \mul/mult_6/U641  ( .A0(n687), .A1(sig_B[7]), .B0(n518), .B1(
        sig_B[6]), .C0(\mul/mult_6/n50 ), .C1(sig_B[5]), .Y(\mul/mult_6/n1147 ) );
  AOI222XL \mul/mult_6/U638  ( .A0(n687), .A1(sig_B[8]), .B0(n518), .B1(
        sig_B[7]), .C0(\mul/mult_6/n50 ), .C1(sig_B[6]), .Y(\mul/mult_6/n1146 ) );
  OAI21X1 \mul/mult_6/U933  ( .A0(n591), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1342 ), .Y(\mul/mult_6/n1316 ) );
  ADDHX1 \mul/mult_6/U269  ( .A(\mul/mult_6/n782 ), .B(\mul/mult_6/n406 ), 
        .CO(\mul/mult_6/n396 ), .S(\mul/mult_6/n397 ) );
  AOI222XL \mul/mult_6/U561  ( .A0(n689), .A1(sig_B[6]), .B0(n690), .B1(
        sig_B[5]), .C0(\mul/mult_6/n60 ), .C1(sig_B[4]), .Y(\mul/mult_6/n1096 ) );
  OAI21X1 \mul/mult_6/U782  ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1243 ), .Y(\mul/mult_6/n1217 ) );
  AOI222XL \mul/mult_6/U555  ( .A0(n689), .A1(sig_B[8]), .B0(n690), .B1(
        sig_B[7]), .C0(\mul/mult_6/n60 ), .C1(sig_B[6]), .Y(\mul/mult_6/n1094 ) );
  OAI21X1 \mul/mult_6/U776  ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1241 ), .Y(\mul/mult_6/n1215 ) );
  OAI21X1 \mul/mult_6/U919  ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1338 ), .Y(\mul/mult_6/n1312 ) );
  ADDFX1 \mul/mult_6/U233  ( .A(n669), .B(n668), .CI(sig_B[5]), .CO(
        \mul/mult_6/n298 ), .S(\mul/mult_6/n299 ) );
  ADDFX1 \mul/mult_6/U210  ( .A(n666), .B(sig_B[9]), .CI(sig_B[11]), .CO(
        \mul/mult_6/n240 ), .S(\mul/mult_6/n241 ) );
  ADDFX1 \mul/mult_6/U193  ( .A(n664), .B(sig_B[15]), .CI(sig_B[17]), .CO(
        \mul/mult_6/n200 ), .S(\mul/mult_6/n201 ) );
  OAI21X1 \mul/mult_6/U1259  ( .A0(\mul/mult_6/n683 ), .A1(\mul/mult_6/n687 ), 
        .B0(\mul/mult_6/n684 ), .Y(\mul/mult_6/n682 ) );
  AND3X6 \mul/mult_6/U1088  ( .A(\mul/mult_6/n1442 ), .B(\mul/mult_6/n1450 ), 
        .C(\mul/mult_6/n1458 ), .Y(\mul/mult_6/n20 ) );
  OAI21X1 \mul/mult_6/U1182  ( .A0(\mul/mult_6/n630 ), .A1(\mul/mult_6/n636 ), 
        .B0(\mul/mult_6/n631 ), .Y(\mul/mult_6/n629 ) );
  NAND2X2 \mul/mult_6/U1256  ( .A(\mul/mult_6/n689 ), .B(\mul/mult_6/n681 ), 
        .Y(\mul/mult_6/n679 ) );
  OAI21X1 \mul/mult_6/U1296  ( .A0(\mul/mult_6/n705 ), .A1(\mul/mult_6/n707 ), 
        .B0(\mul/mult_6/n706 ), .Y(\mul/mult_6/n704 ) );
  ADDFX1 \sub/sub_17/U7  ( .A(\sub/sub_17/n15 ), .B(exp_C[2]), .CI(
        \sub/sub_17/n7 ), .CO(\sub/sub_17/n6 ), .S(\sub/N16 ) );
  ADDFX1 \sub/r301/U7  ( .A(exp_P[2]), .B(n1061), .CI(\sub/r301/n7 ), .CO(
        \sub/r301/n6 ), .S(\sub/N7 ) );
  OAI21X1 \mul/mult_6/U496  ( .A0(n678), .A1(\mul/mult_6/n68 ), .B0(n586), .Y(
        \mul/mult_6/n1024 ) );
  OAI21X1 \mul/mult_6/U492  ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n68 ), 
        .B0(n610), .Y(\mul/mult_6/n1023 ) );
  OAI21X1 \mul/mult_6/U489  ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1048 ), .Y(\mul/mult_6/n1022 ) );
  ADDFX1 \sub/r301/U6  ( .A(exp_P[3]), .B(n1049), .CI(\sub/r301/n6 ), .CO(
        \sub/r301/n5 ), .S(\sub/N8 ) );
  ADDFX1 \sub/sub_17/U6  ( .A(\sub/sub_17/n14 ), .B(exp_C[3]), .CI(
        \sub/sub_17/n6 ), .CO(\sub/sub_17/n5 ), .S(\sub/N17 ) );
  AOI21X1 \mul/mult_6/U1279  ( .A0(\mul/mult_6/n698 ), .A1(\mul/mult_6/n729 ), 
        .B0(\mul/mult_6/n695 ), .Y(\mul/mult_6/n693 ) );
  ADDFX1 \sub/sub_17/U5  ( .A(n1046), .B(exp_C[4]), .CI(\sub/sub_17/n5 ), .CO(
        \sub/sub_17/n4 ), .S(\sub/N18 ) );
  OAI21X1 \mul/mult_6/U1265  ( .A0(\mul/mult_6/n688 ), .A1(\mul/mult_6/n686 ), 
        .B0(\mul/mult_6/n687 ), .Y(\mul/mult_6/n685 ) );
  OAI21X1 \mul/mult_6/U815  ( .A0(n545), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1254 ), .Y(\mul/mult_6/n1228 ) );
  ADDFX1 \sub/r301/U5  ( .A(exp_P[4]), .B(\sub/r301/n13 ), .CI(\sub/r301/n5 ), 
        .CO(\sub/r301/n4 ), .S(\sub/N9 ) );
  ADDFX1 \sub/r301/U4  ( .A(exp_P[5]), .B(n1029), .CI(\sub/r301/n4 ), .CO(
        \sub/r301/n3 ), .S(\sub/N10 ) );
  ADDFX1 \sub/sub_17/U4  ( .A(n1047), .B(exp_C[5]), .CI(\sub/sub_17/n4 ), .CO(
        \sub/sub_17/n3 ), .S(\sub/N19 ) );
  ADDHX1 \mul/mult_6/U305  ( .A(\mul/mult_6/n488 ), .B(\mul/mult_6/n891 ), 
        .CO(\mul/mult_6/n484 ), .S(\mul/mult_6/n485 ) );
  ADDFX1 \mul/mult_6/U185  ( .A(n670), .B(\mul/mult_6/n186 ), .CI(n541), .CO(
        \mul/mult_6/n183 ), .S(\mul/mult_6/n184 ) );
  OAI21X1 \mul/mult_6/U889  ( .A0(n544), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1303 ), .Y(\mul/mult_6/n1277 ) );
  OAI21X1 \mul/mult_6/U803  ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1250 ), .Y(\mul/mult_6/n1224 ) );
  OAI21X1 \mul/mult_6/U729  ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1201 ), .Y(\mul/mult_6/n1175 ) );
  OAI21X1 \mul/mult_6/U963  ( .A0(n542), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1352 ), .Y(\mul/mult_6/n1326 ) );
  OAI21X1 \mul/mult_6/U856  ( .A0(n569), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1292 ), .Y(\mul/mult_6/n1266 ) );
  OAI21X1 \mul/mult_6/U945  ( .A0(n570), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1346 ), .Y(\mul/mult_6/n1320 ) );
  OAI21X1 \mul/mult_6/U806  ( .A0(n544), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1251 ), .Y(\mul/mult_6/n1225 ) );
  OAI21X1 \mul/mult_6/U978  ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1357 ), .Y(\mul/mult_6/n1331 ) );
  OAI21X1 \mul/mult_6/U880  ( .A0(n542), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1300 ), .Y(\mul/mult_6/n1274 ) );
  ADDHX1 \mul/mult_6/U299  ( .A(\mul/mult_6/n476 ), .B(\mul/mult_6/n864 ), 
        .CO(\mul/mult_6/n471 ), .S(\mul/mult_6/n472 ) );
  OAI21X1 \mul/mult_6/U883  ( .A0(n543), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1301 ), .Y(\mul/mult_6/n1275 ) );
  OAI21X1 \mul/mult_6/U886  ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1302 ), .Y(\mul/mult_6/n1276 ) );
  ADDFX1 \sub/r301/U3  ( .A(exp_P[6]), .B(n1032), .CI(\sub/r301/n3 ), .CO(
        \sub/r301/n2 ), .S(\sub/N11 ) );
  OAI21X1 \mul/mult_6/U812  ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1253 ), .Y(\mul/mult_6/n1227 ) );
  ADDFX1 \sub/sub_17/U3  ( .A(n1031), .B(exp_C[6]), .CI(\sub/sub_17/n3 ), .CO(
        \sub/sub_17/n2 ), .S(\sub/N20 ) );
  OAI21X1 \mul/mult_6/U951  ( .A0(n571), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1348 ), .Y(\mul/mult_6/n1322 ) );
  OAI21X1 \mul/mult_6/U862  ( .A0(n570), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1294 ), .Y(\mul/mult_6/n1268 ) );
  OAI21X1 \mul/mult_6/U868  ( .A0(n571), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1296 ), .Y(\mul/mult_6/n1270 ) );
  OAI21X1 \mul/mult_6/U939  ( .A0(n569), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1344 ), .Y(\mul/mult_6/n1318 ) );
  OAI21X1 \mul/mult_6/U957  ( .A0(n572), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1350 ), .Y(\mul/mult_6/n1324 ) );
  ADDHX1 \mul/mult_6/U280  ( .A(\mul/mult_6/n809 ), .B(\mul/mult_6/n432 ), 
        .CO(\mul/mult_6/n424 ), .S(\mul/mult_6/n425 ) );
  ADDFX1 \mul/mult_6/U253  ( .A(sig_B[0]), .B(n606), .CI(\mul/mult_6/n364 ), 
        .CO(\mul/mult_6/n353 ), .S(\mul/mult_6/n354 ) );
  ADDHX1 \mul/mult_6/U297  ( .A(\mul/mult_6/n863 ), .B(\mul/mult_6/n471 ), 
        .CO(\mul/mult_6/n466 ), .S(\mul/mult_6/n467 ) );
  ADDFX1 \mul/mult_6/U245  ( .A(sig_A[2]), .B(sig_B[2]), .CI(n607), .CO(
        \mul/mult_6/n331 ), .S(\mul/mult_6/n332 ) );
  ADDFX1 \mul/mult_6/U241  ( .A(sig_A[2]), .B(sig_B[3]), .CI(n628), .CO(
        \mul/mult_6/n320 ), .S(\mul/mult_6/n321 ) );
  OAI21X1 \mul/mult_6/U865  ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1295 ), .Y(\mul/mult_6/n1269 ) );
  OAI21X1 \mul/mult_6/U927  ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1340 ), .Y(\mul/mult_6/n1314 ) );
  ADDFX1 \mul/mult_6/U237  ( .A(sig_A[2]), .B(sig_B[4]), .CI(\mul/mult_6/n320 ), .CO(\mul/mult_6/n309 ), .S(\mul/mult_6/n310 ) );
  OAI21X1 \mul/mult_6/U853  ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1291 ), .Y(\mul/mult_6/n1265 ) );
  ADDHX1 \mul/mult_6/U173  ( .A(\mul/mult_6/n173 ), .B(\mul/mult_6/n944 ), 
        .CO(\mul/mult_6/n172 ), .S(sig_P[2]) );
  OAI21X1 \mul/mult_6/U794  ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1247 ), .Y(\mul/mult_6/n1221 ) );
  OAI21X1 \mul/mult_6/U948  ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1347 ), .Y(\mul/mult_6/n1321 ) );
  OAI21X1 \mul/mult_6/U923  ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1339 ), .Y(\mul/mult_6/n1313 ) );
  OAI21X1 \mul/mult_6/U930  ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1341 ), .Y(\mul/mult_6/n1315 ) );
  OAI21X1 \mul/mult_6/U942  ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1345 ), .Y(\mul/mult_6/n1319 ) );
  OAI21X1 \mul/mult_6/U859  ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1293 ), .Y(\mul/mult_6/n1267 ) );
  OAI21X1 \mul/mult_6/U871  ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1297 ), .Y(\mul/mult_6/n1271 ) );
  OAI21X1 \mul/mult_6/U877  ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1299 ), .Y(\mul/mult_6/n1273 ) );
  OAI21X1 \mul/mult_6/U954  ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1349 ), .Y(\mul/mult_6/n1323 ) );
  OAI21X1 \mul/mult_6/U936  ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1343 ), .Y(\mul/mult_6/n1317 ) );
  OAI21X1 \mul/mult_6/U960  ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1351 ), .Y(\mul/mult_6/n1325 ) );
  MXI2XL \align/sra_11/U432  ( .A(\align/sra_11/n563 ), .B(\align/sra_11/n564 ), .S0(n718), .Y(\align/sra_11/n562 ) );
  MXI2XL \align/sra_11/U615  ( .A(\align/sra_11/n534 ), .B(\align/sra_11/n535 ), .S0(n717), .Y(\align/sra_11/n533 ) );
  MXI2XL \align/sra_11/U501  ( .A(\align/sra_11/n633 ), .B(\align/sra_11/n558 ), .S0(n717), .Y(\align/sra_11/n632 ) );
  MXI2X2 \align/sra_10/U254  ( .A(\align/sra_10/n300 ), .B(\align/sra_10/n301 ), .S0(n507), .Y(\align/sra_10/n246 ) );
  MXI2X2 \align/sra_10/U201  ( .A(\align/sra_10/n249 ), .B(n706), .S0(
        \align/sra_11/SH[1] ), .Y(\align/sra_10/n199 ) );
  MXI2X2 \align/sra_10/U117  ( .A(\align/sra_10/n133 ), .B(\align/sra_10/n141 ), .S0(n705), .Y(\align/sra_10/n83 ) );
  MXI2X2 \align/sra_10/U82  ( .A(\align/sra_10/n68 ), .B(\align/sra_10/n100 ), 
        .S0(n717), .Y(\align/sra_10/n18 ) );
  AOI21X2 \sigadd/add_9/U329  ( .A0(\sigadd/add_9/n242 ), .A1(n553), .B0(
        \sigadd/add_9/n239 ), .Y(\sigadd/add_9/n237 ) );
  AOI21X4 \sigadd/add_9/U315  ( .A0(\sigadd/add_9/n234 ), .A1(n552), .B0(
        \sigadd/add_9/n231 ), .Y(\sigadd/add_9/n229 ) );
  OAI21X4 \sigadd/add_9/U309  ( .A0(\sigadd/add_9/n229 ), .A1(
        \sigadd/add_9/n227 ), .B0(\sigadd/add_9/n228 ), .Y(\sigadd/add_9/n226 ) );
  AOI21X4 \sigadd/add_9/U301  ( .A0(\sigadd/add_9/n226 ), .A1(n551), .B0(
        \sigadd/add_9/n223 ), .Y(\sigadd/add_9/n221 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U6  ( .A(n559), .B(\sigadd/sub_add_11_b0/n6 ), 
        .CO(\sigadd/sub_add_11_b0/n5 ), .S(\sigadd/N46 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U5  ( .A(n566), .B(\sigadd/sub_add_11_b0/n5 ), 
        .CO(\sigadd/sub_add_11_b0/n4 ), .S(\sigadd/N47 ) );
  MXI2XL \normal/srl_15/U293  ( .A(\normal/srl_15/A[1] ), .B(add_out[17]), 
        .S0(n703), .Y(\normal/srl_15/n200 ) );
  MXI2XL \normal/srl_15/U294  ( .A(\sigadd/sig[0] ), .B(add_out[16]), .S0(n703), .Y(\normal/srl_15/n199 ) );
  MXI2XL \normal/sll_15/U236  ( .A(add_out[45]), .B(\normal/srl_15/A[29] ), 
        .S0(n714), .Y(\normal/sll_15/n234 ) );
  MXI2XL \normal/sll_15/U235  ( .A(add_out[46]), .B(add_out[30]), .S0(n703), 
        .Y(\normal/sll_15/n235 ) );
  MXI2XL \normal/srl_15/U242  ( .A(\normal/srl_15/n201 ), .B(
        \normal/srl_15/n203 ), .S0(n715), .Y(\normal/srl_15/n151 ) );
  MXI2XL \normal/srl_15/U243  ( .A(\normal/srl_15/n200 ), .B(
        \normal/srl_15/n202 ), .S0(n715), .Y(\normal/srl_15/n150 ) );
  MXI2XL \normal/srl_15/U241  ( .A(\normal/srl_15/n202 ), .B(
        \normal/srl_15/n204 ), .S0(n715), .Y(\normal/srl_15/n152 ) );
  MXI2XL \normal/srl_15/U237  ( .A(\normal/srl_15/n206 ), .B(
        \normal/srl_15/n208 ), .S0(n715), .Y(\normal/srl_15/n156 ) );
  MXI2XL \normal/srl_15/U238  ( .A(\normal/srl_15/n205 ), .B(
        \normal/srl_15/n207 ), .S0(n715), .Y(\normal/srl_15/n155 ) );
  MXI2XL \normal/srl_15/U239  ( .A(\normal/srl_15/n204 ), .B(
        \normal/srl_15/n206 ), .S0(n715), .Y(\normal/srl_15/n154 ) );
  MXI2XL \normal/srl_15/U240  ( .A(\normal/srl_15/n203 ), .B(
        \normal/srl_15/n205 ), .S0(n715), .Y(\normal/srl_15/n153 ) );
  MXI2XL \normal/srl_15/U244  ( .A(\normal/srl_15/n199 ), .B(
        \normal/srl_15/n201 ), .S0(n715), .Y(\normal/srl_15/n149 ) );
  MXI2XL \normal/srl_15/U191  ( .A(\normal/srl_15/n152 ), .B(
        \normal/srl_15/n184 ), .S0(n504), .Y(\normal/srl_15/n102 ) );
  NAND2X2 \ctrl/add_1_root_add_16_2/U61  ( .A(n520), .B(n534), .Y(
        \ctrl/add_1_root_add_16_2/n48 ) );
  XNOR2X1 \ctrl/sub_0_root_add_0_root_sub_16/U47  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[0] ), .B(n711), .Y(\ctrl/N27 ) );
  XNOR2X1 \ctrl/add_1_root_add_16_2/U69  ( .A(n702), .B(
        \ctrl/add_1_root_add_16_2/n6 ), .Y(\ctrl/N11 ) );
  AND3X6 \mul/mult_6/U1067  ( .A(\mul/mult_6/n1439 ), .B(\mul/mult_6/n1447 ), 
        .C(\mul/mult_6/n1455 ), .Y(\mul/mult_6/n50 ) );
  XOR2X1 \mul/mult_6/U1295  ( .A(\mul/mult_6/n572 ), .B(\mul/mult_6/n707 ), 
        .Y(\mul/mult_6/n1411 ) );
  AND3X6 \mul/mult_6/U1095  ( .A(\mul/mult_6/n1451 ), .B(\mul/mult_6/n1459 ), 
        .C(\mul/mult_6/n1443 ), .Y(\mul/mult_6/n9 ) );
  NAND2X2 \mul/mult_6/U1140  ( .A(\mul/mult_6/n613 ), .B(\mul/mult_6/n601 ), 
        .Y(\mul/mult_6/n599 ) );
  NAND2X2 \mul/mult_6/U1179  ( .A(\mul/mult_6/n640 ), .B(\mul/mult_6/n628 ), 
        .Y(\mul/mult_6/n626 ) );
  AOI21X1 \mul/mult_6/U1180  ( .A0(\mul/mult_6/n628 ), .A1(\mul/mult_6/n643 ), 
        .B0(\mul/mult_6/n629 ), .Y(\mul/mult_6/n627 ) );
  NAND2X2 \mul/mult_6/U1114  ( .A(\mul/mult_6/n589 ), .B(n592), .Y(
        \mul/mult_6/n582 ) );
  NOR2X2 \mul/mult_6/U1177  ( .A(\mul/mult_6/n652 ), .B(\mul/mult_6/n626 ), 
        .Y(\mul/mult_6/n624 ) );
  XOR2X1 \expadd/add_0_root_sub_0_root_sub_8/U2  ( .A(
        \expadd/add_0_root_sub_0_root_sub_8/B[7] ), .B(exp_B[7]), .Y(
        \expadd/add_0_root_sub_0_root_sub_8/n1 ) );
  OAI21X1 \mul/mult_6/U486  ( .A0(n546), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1047 ), .Y(\mul/mult_6/n1021 ) );
  AOI21X1 \mul/mult_6/U1198  ( .A0(\mul/mult_6/n655 ), .A1(\mul/mult_6/n640 ), 
        .B0(\mul/mult_6/n643 ), .Y(\mul/mult_6/n639 ) );
  NOR2X2 \mul/mult_6/U1106  ( .A(\mul/mult_6/n581 ), .B(sig_B[22]), .Y(
        \mul/mult_6/n576 ) );
  XOR2X1 \mul/mult_6/U485  ( .A(\mul/mult_6/n1021 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n781 ) );
  XOR2X1 \mul/mult_6/U495  ( .A(\mul/mult_6/n1024 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n784 ) );
  OAI21X1 \mul/mult_6/U981  ( .A0(n545), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1358 ), .Y(\mul/mult_6/n1332 ) );
  XOR2X1 \mul/mult_6/U488  ( .A(\mul/mult_6/n1022 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n782 ) );
  XOR2X1 \mul/mult_6/U491  ( .A(\mul/mult_6/n1023 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n783 ) );
  XOR2XL \mul/mult_6/U989  ( .A(\mul/mult_6/n1335 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n945 ) );
  OAI21X1 \mul/mult_6/U566  ( .A0(n545), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1098 ), .Y(\mul/mult_6/n1072 ) );
  XOR2XL \mul/mult_6/U983  ( .A(\mul/mult_6/n1333 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n943 ) );
  OAI21X1 \mul/mult_6/U587  ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1130 ), .Y(\mul/mult_6/n1104 ) );
  OAI21X1 \mul/mult_6/U421  ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1026 ), .Y(\mul/mult_6/n1000 ) );
  ADDHX1 \mul/mult_6/U277  ( .A(sig_A[20]), .B(\mul/mult_6/n784 ), .CO(
        \mul/mult_6/n416 ), .S(\mul/mult_6/n417 ) );
  XOR2X1 \mul/mult_6/U814  ( .A(\mul/mult_6/n1228 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n888 ) );
  OAI21X1 \mul/mult_6/U504  ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1078 ), .Y(\mul/mult_6/n1052 ) );
  XOR2X1 \mul/mult_6/U482  ( .A(\mul/mult_6/n1020 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n780 ) );
  XOR2X1 \mul/mult_6/U503  ( .A(\mul/mult_6/n1052 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n787 ) );
  XOR2X1 \mul/mult_6/U1195  ( .A(\mul/mult_6/n646 ), .B(\mul/mult_6/n561 ), 
        .Y(\mul/mult_6/n1400 ) );
  OAI21X1 \mul/mult_6/U557  ( .A0(n544), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1095 ), .Y(\mul/mult_6/n1069 ) );
  OAI21X1 \mul/mult_6/U966  ( .A0(n543), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1353 ), .Y(\mul/mult_6/n1327 ) );
  OAI21X1 \mul/mult_6/U560  ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1096 ), .Y(\mul/mult_6/n1070 ) );
  OAI21X1 \mul/mult_6/U584  ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n48 ), 
        .B0(n688), .Y(\mul/mult_6/n1103 ) );
  OAI21X1 \mul/mult_6/U563  ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1097 ), .Y(\mul/mult_6/n1071 ) );
  XOR2X1 \mul/mult_6/U420  ( .A(\mul/mult_6/n1000 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n760 ) );
  OAI21X1 \mul/mult_6/U418  ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n68 ), 
        .B0(n694), .Y(\mul/mult_6/n999 ) );
  ADDHX1 \mul/mult_6/U309  ( .A(\mul/mult_6/n494 ), .B(\mul/mult_6/n918 ), 
        .CO(\mul/mult_6/n492 ), .S(\mul/mult_6/n493 ) );
  OAI21X1 \mul/mult_6/U501  ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n58 ), 
        .B0(n691), .Y(\mul/mult_6/n1051 ) );
  ADDHX1 \mul/mult_6/U303  ( .A(\mul/mult_6/n890 ), .B(\mul/mult_6/n484 ), 
        .CO(\mul/mult_6/n480 ), .S(\mul/mult_6/n481 ) );
  ADDHX1 \mul/mult_6/U308  ( .A(\mul/mult_6/n917 ), .B(\mul/mult_6/n492 ), 
        .CO(\mul/mult_6/n490 ), .S(\mul/mult_6/n491 ) );
  XOR2X1 \mul/mult_6/U500  ( .A(\mul/mult_6/n1051 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n786 ) );
  ADDHX1 \mul/mult_6/U174  ( .A(\mul/mult_6/n176 ), .B(\mul/mult_6/n945 ), 
        .CO(\mul/mult_6/n173 ), .S(sig_P[1]) );
  XOR2X1 \mul/mult_6/U434  ( .A(\mul/mult_6/n1004 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n764 ) );
  XOR2X1 \mul/mult_6/U417  ( .A(\mul/mult_6/n999 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n759 ) );
  OAI21X1 \mul/mult_6/U432  ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1029 ), .Y(\mul/mult_6/n1003 ) );
  OAI21X1 \mul/mult_6/U425  ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1027 ), .Y(\mul/mult_6/n1001 ) );
  XOR2X1 \mul/mult_6/U507  ( .A(\mul/mult_6/n1053 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n788 ) );
  XOR2X1 \mul/mult_6/U437  ( .A(\mul/mult_6/n1005 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n765 ) );
  XOR2X1 \mul/mult_6/U511  ( .A(\mul/mult_6/n1054 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n789 ) );
  XOR2X1 \mul/mult_6/U424  ( .A(\mul/mult_6/n1001 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n761 ) );
  ADDFX1 \mul/mult_6/U304  ( .A(\mul/mult_6/n485 ), .B(\mul/mult_6/n915 ), 
        .CI(\mul/mult_6/n486 ), .CO(\mul/mult_6/n482 ), .S(\mul/mult_6/n483 )
         );
  XOR2X1 \mul/mult_6/U514  ( .A(\mul/mult_6/n1055 ), .B(sig_A[17]), .Y(
        \mul/mult_6/n790 ) );
  ADDFX1 \mul/mult_6/U168  ( .A(\mul/mult_6/n939 ), .B(\mul/mult_6/n483 ), 
        .CI(\mul/mult_6/n168 ), .CO(\mul/mult_6/n167 ), .S(sig_P[7]) );
  ADDFX1 \mul/mult_6/U167  ( .A(\mul/mult_6/n479 ), .B(\mul/mult_6/n482 ), 
        .CI(\mul/mult_6/n167 ), .CO(\mul/mult_6/n166 ), .S(sig_P[8]) );
  MXI2XL \align/sra_11/U474  ( .A(\align/sra_11/n518 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n517 ) );
  MXI2XL \align/sra_11/U446  ( .A(\align/sra_11/n516 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n515 ) );
  MXI2X1 \align/sra_11/U704  ( .A(\align/sra_11/n718 ), .B(\align/sra_11/n587 ), .S0(n719), .Y(\align/sra_11/n715 ) );
  MXI2X1 \align/sra_11/U697  ( .A(\align/sra_11/n697 ), .B(\align/sra_11/n583 ), .S0(n719), .Y(\align/sra_11/n694 ) );
  MXI2X1 \align/sra_11/U431  ( .A(\align/sra_11/n567 ), .B(\align/sra_11/n568 ), .S0(n718), .Y(\align/sra_11/n566 ) );
  MXI2X1 \align/sra_11/U691  ( .A(\align/sra_11/n684 ), .B(\align/sra_11/n567 ), .S0(n719), .Y(\align/sra_11/n682 ) );
  MXI2X1 \align/sra_11/U430  ( .A(\align/sra_11/n583 ), .B(\align/sra_11/n584 ), .S0(n718), .Y(\align/sra_11/n582 ) );
  MXI2X1 \align/sra_11/U428  ( .A(\align/sra_11/n591 ), .B(\align/sra_11/n592 ), .S0(n718), .Y(\align/sra_11/n590 ) );
  MXI2X1 \align/sra_11/U429  ( .A(\align/sra_11/n587 ), .B(\align/sra_11/n588 ), .S0(n718), .Y(\align/sra_11/n586 ) );
  MXI2X1 \align/sra_11/U685  ( .A(\align/sra_11/n672 ), .B(\align/sra_11/n563 ), .S0(n719), .Y(\align/sra_11/n670 ) );
  MXI2XL \align/sra_11/U443  ( .A(\align/sra_11/n526 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n525 ) );
  MXI2XL \align/sra_11/U442  ( .A(\align/sra_11/n528 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n527 ) );
  MXI2XL \align/sra_11/U473  ( .A(\align/sra_11/n520 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n519 ) );
  MXI2XL \align/sra_11/U444  ( .A(\align/sra_11/n524 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n523 ) );
  MXI2XL \align/sra_11/U441  ( .A(\align/sra_11/n467 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n529 ) );
  MXI2XL \align/sra_11/U633  ( .A(\align/sra_11/n570 ), .B(\align/sra_11/n556 ), .S0(n515), .Y(\align/sra_11/n569 ) );
  MXI2XL \align/sra_11/U445  ( .A(\align/sra_11/n522 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n521 ) );
  MXI2XL \align/sra_11/U728  ( .A(\align/sra_11/n754 ), .B(\align/sra_11/n757 ), .S0(n515), .Y(\align/sra_11/n753 ) );
  ADDFHX2 \mul/mult_6/U148  ( .A(\mul/mult_6/n313 ), .B(\mul/mult_6/n323 ), 
        .CI(\mul/mult_6/n148 ), .CO(\mul/mult_6/n147 ), .S(sig_P[27]) );
  MXI2X2 \align/sra_10/U252  ( .A(\align/sra_10/n302 ), .B(\align/sra_10/n303 ), .S0(n507), .Y(\align/sra_10/n248 ) );
  MXI2X2 \align/sra_10/U256  ( .A(\align/sra_10/n298 ), .B(\align/sra_10/n299 ), .S0(n507), .Y(\align/sra_10/n244 ) );
  MXI2X1 \align/sra_10/U121  ( .A(\align/sra_10/n129 ), .B(\align/sra_10/n137 ), .S0(n705), .Y(\align/sra_10/n79 ) );
  MXI2X1 \align/sra_10/U128  ( .A(\align/sra_10/n122 ), .B(\align/sra_10/n130 ), .S0(n506), .Y(\align/sra_10/n72 ) );
  MXI2X1 \align/sra_10/U127  ( .A(\align/sra_10/n123 ), .B(\align/sra_10/n131 ), .S0(n506), .Y(\align/sra_10/n73 ) );
  MXI2X1 \align/sra_10/U122  ( .A(\align/sra_10/n128 ), .B(\align/sra_10/n136 ), .S0(n705), .Y(\align/sra_10/n78 ) );
  MXI2X1 \align/sra_10/U120  ( .A(\align/sra_10/n130 ), .B(\align/sra_10/n138 ), .S0(n705), .Y(\align/sra_10/n80 ) );
  MXI2X1 \align/sra_10/U129  ( .A(\align/sra_10/n121 ), .B(\align/sra_10/n129 ), .S0(n506), .Y(\align/sra_10/n71 ) );
  MXI2X1 \align/sra_10/U124  ( .A(\align/sra_10/n126 ), .B(\align/sra_10/n134 ), .S0(n705), .Y(\align/sra_10/n76 ) );
  MXI2X1 \align/sra_10/U126  ( .A(\align/sra_10/n124 ), .B(\align/sra_10/n132 ), .S0(n506), .Y(\align/sra_10/n74 ) );
  MXI2X1 \align/sra_10/U119  ( .A(\align/sra_10/n131 ), .B(\align/sra_10/n139 ), .S0(n705), .Y(\align/sra_10/n81 ) );
  MXI2X1 \align/sra_10/U123  ( .A(\align/sra_10/n127 ), .B(\align/sra_10/n135 ), .S0(n705), .Y(\align/sra_10/n77 ) );
  MXI2X1 \align/sra_10/U125  ( .A(\align/sra_10/n125 ), .B(\align/sra_10/n133 ), .S0(n705), .Y(\align/sra_10/n75 ) );
  MXI2X1 \align/sra_10/U118  ( .A(\align/sra_10/n132 ), .B(\align/sra_10/n140 ), .S0(n705), .Y(\align/sra_10/n82 ) );
  NAND2X2 \sigadd/add_9/U209  ( .A(ali_P[20]), .B(ali_C[20]), .Y(
        \sigadd/add_9/n169 ) );
  NAND2X2 \sigadd/add_9/U167  ( .A(ali_P[26]), .B(ali_C[26]), .Y(
        \sigadd/add_9/n145 ) );
  NAND2X2 \sigadd/add_9/U139  ( .A(ali_P[30]), .B(ali_C[30]), .Y(
        \sigadd/add_9/n129 ) );
  NAND2X2 \sigadd/add_9/U181  ( .A(ali_P[24]), .B(ali_C[24]), .Y(
        \sigadd/add_9/n153 ) );
  NAND2X2 \sigadd/add_9/U47  ( .A(ali_P[43]), .B(ali_C[43]), .Y(
        \sigadd/add_9/n76 ) );
  NAND2X2 \sigadd/add_9/U19  ( .A(ali_P[47]), .B(ali_C[47]), .Y(
        \sigadd/add_9/n60 ) );
  NAND2X2 \sigadd/add_9/U195  ( .A(ali_P[22]), .B(ali_C[22]), .Y(
        \sigadd/add_9/n161 ) );
  NAND2X2 \sigadd/add_9/U257  ( .A(ali_P[13]), .B(ali_C[13]), .Y(
        \sigadd/add_9/n196 ) );
  NAND2X2 \sigadd/add_9/U89  ( .A(ali_P[37]), .B(ali_C[37]), .Y(
        \sigadd/add_9/n100 ) );
  NAND2X2 \sigadd/add_9/U33  ( .A(ali_P[45]), .B(ali_C[45]), .Y(
        \sigadd/add_9/n68 ) );
  NAND2X2 \sigadd/add_9/U251  ( .A(ali_P[14]), .B(ali_C[14]), .Y(
        \sigadd/add_9/n193 ) );
  NAND2X2 \sigadd/add_9/U61  ( .A(ali_P[41]), .B(ali_C[41]), .Y(
        \sigadd/add_9/n84 ) );
  NAND2X2 \sigadd/add_9/U75  ( .A(ali_P[39]), .B(ali_C[39]), .Y(
        \sigadd/add_9/n92 ) );
  NAND2X2 \sigadd/add_9/U237  ( .A(ali_P[16]), .B(ali_C[16]), .Y(
        \sigadd/add_9/n185 ) );
  NAND2X2 \sigadd/add_9/U153  ( .A(ali_P[28]), .B(ali_C[28]), .Y(
        \sigadd/add_9/n137 ) );
  NAND2XL \sigadd/add_9/U304  ( .A(n551), .B(\sigadd/add_9/n225 ), .Y(
        \sigadd/add_9/n44 ) );
  NAND2XL \sigadd/add_9/U290  ( .A(n550), .B(\sigadd/add_9/n217 ), .Y(
        \sigadd/add_9/n42 ) );
  NAND2XL \sigadd/add_9/U262  ( .A(n548), .B(\sigadd/add_9/n201 ), .Y(
        \sigadd/add_9/n38 ) );
  NAND2XL \sigadd/add_9/U276  ( .A(n549), .B(\sigadd/add_9/n209 ), .Y(
        \sigadd/add_9/n40 ) );
  NAND2XL \sigadd/add_9/U332  ( .A(n553), .B(\sigadd/add_9/n241 ), .Y(
        \sigadd/add_9/n48 ) );
  NAND2XL \sigadd/add_9/U318  ( .A(n552), .B(\sigadd/add_9/n233 ), .Y(
        \sigadd/add_9/n46 ) );
  NAND2XL \sigadd/add_9/U324  ( .A(\sigadd/add_9/n293 ), .B(
        \sigadd/add_9/n236 ), .Y(\sigadd/add_9/n47 ) );
  NAND2XL \sigadd/add_9/U296  ( .A(\sigadd/add_9/n289 ), .B(
        \sigadd/add_9/n220 ), .Y(\sigadd/add_9/n43 ) );
  NAND2XL \sigadd/add_9/U310  ( .A(\sigadd/add_9/n291 ), .B(
        \sigadd/add_9/n228 ), .Y(\sigadd/add_9/n45 ) );
  NAND2XL \sigadd/add_9/U254  ( .A(\sigadd/add_9/n283 ), .B(
        \sigadd/add_9/n196 ), .Y(\sigadd/add_9/n37 ) );
  NAND2XL \sigadd/add_9/U30  ( .A(\sigadd/add_9/n251 ), .B(\sigadd/add_9/n68 ), 
        .Y(\sigadd/add_9/n5 ) );
  NAND2XL \sigadd/add_9/U240  ( .A(\sigadd/add_9/n281 ), .B(
        \sigadd/add_9/n188 ), .Y(\sigadd/add_9/n35 ) );
  NAND2XL \sigadd/add_9/U268  ( .A(\sigadd/add_9/n285 ), .B(
        \sigadd/add_9/n204 ), .Y(\sigadd/add_9/n39 ) );
  NAND2XL \sigadd/add_9/U282  ( .A(\sigadd/add_9/n287 ), .B(
        \sigadd/add_9/n212 ), .Y(\sigadd/add_9/n41 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U16  ( .A(n584), .B(\sigadd/sub_add_11_b0/n16 ), 
        .CO(\sigadd/sub_add_11_b0/n15 ), .S(\sigadd/N36 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U15  ( .A(n590), .B(\sigadd/sub_add_11_b0/n15 ), 
        .CO(\sigadd/sub_add_11_b0/n14 ), .S(\sigadd/N37 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U14  ( .A(n583), .B(\sigadd/sub_add_11_b0/n14 ), 
        .CO(\sigadd/sub_add_11_b0/n13 ), .S(\sigadd/N38 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U13  ( .A(n589), .B(\sigadd/sub_add_11_b0/n13 ), 
        .CO(\sigadd/sub_add_11_b0/n12 ), .S(\sigadd/N39 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U7  ( .A(n567), .B(\sigadd/sub_add_11_b0/n7 ), 
        .CO(\sigadd/sub_add_11_b0/n6 ), .S(\sigadd/N45 ) );
  MXI2XL \normal/srl_15/U236  ( .A(\normal/srl_15/n207 ), .B(
        \normal/srl_15/n209 ), .S0(n715), .Y(\normal/srl_15/n157 ) );
  MXI2XL \normal/srl_15/U193  ( .A(\normal/srl_15/n150 ), .B(
        \normal/srl_15/n182 ), .S0(n504), .Y(\normal/srl_15/n100 ) );
  NAND2X2 \ctrl/add_1_root_add_16_2/U18  ( .A(n504), .B(mux_out[5]), .Y(
        \ctrl/add_1_root_add_16_2/n19 ) );
  MXI2XL \normal/srl_15/U194  ( .A(\normal/srl_15/n149 ), .B(
        \normal/srl_15/n181 ), .S0(n504), .Y(\normal/srl_15/n99 ) );
  MXI2XL \normal/srl_15/U192  ( .A(\normal/srl_15/n151 ), .B(
        \normal/srl_15/n183 ), .S0(n504), .Y(\normal/srl_15/n101 ) );
  MXI2X1 \normal/sll_15/U7  ( .A(\normal/sll_15/n41 ), .B(\normal/sll_15/n40 ), 
        .S0(n503), .Y(\normal/N88 ) );
  NAND2X4 \round/r298/U93  ( .A(norm_out[12]), .B(norm_out[13]), .Y(
        \round/r298/n76 ) );
  NAND2X4 \round/r298/U65  ( .A(norm_out[17]), .B(norm_out[16]), .Y(
        \round/r298/n52 ) );
  NOR2X2 \ctrl/add_1_root_add_16_2/U13  ( .A(\ctrl/add_1_root_add_16_2/n23 ), 
        .B(\ctrl/add_1_root_add_16_2/n18 ), .Y(\ctrl/add_1_root_add_16_2/n16 )
         );
  NOR2X4 \round/r298/U140  ( .A(n522), .B(\round/r298/n117 ), .Y(
        \round/r298/n116 ) );
  NAND2X4 \round/r298/U136  ( .A(\round/r298/n116 ), .B(norm_out[5]), .Y(
        \round/r298/n113 ) );
  XOR2X1 \ctrl/add_1_root_add_16_2/U31  ( .A(\ctrl/add_1_root_add_16_2/n38 ), 
        .B(\ctrl/add_1_root_add_16_2/n3 ), .Y(\ctrl/N14 ) );
  XOR2X1 \ctrl/add_1_root_add_16_2/U53  ( .A(\ctrl/add_1_root_add_16_2/n58 ), 
        .B(\ctrl/add_1_root_add_16_2/n5 ), .Y(\ctrl/N12 ) );
  NAND2X2 \ctrl/sub_0_root_add_0_root_sub_16/U46  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[1] ), .B(n710), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n34 ) );
  NAND2X2 \ctrl/sub_0_root_add_0_root_sub_16/U40  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[2] ), .B(n712), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n31 ) );
  OAI21X4 \ctrl/sub_0_root_add_0_root_sub_16/U28  ( .A0(
        \ctrl/sub_0_root_add_0_root_sub_16/n27 ), .A1(
        \ctrl/sub_0_root_add_0_root_sub_16/n25 ), .B0(
        \ctrl/sub_0_root_add_0_root_sub_16/n26 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n24 ) );
  OAI21X2 \ctrl/sub_0_root_add_0_root_sub_16/U10  ( .A0(
        \ctrl/sub_0_root_add_0_root_sub_16/n19 ), .A1(
        \ctrl/sub_0_root_add_0_root_sub_16/n8 ), .B0(
        \ctrl/sub_0_root_add_0_root_sub_16/n14 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n12 ) );
  OAI21X1 \mul/mult_6/U1290  ( .A0(\mul/mult_6/n702 ), .A1(\mul/mult_6/n706 ), 
        .B0(\mul/mult_6/n703 ), .Y(\mul/mult_6/n701 ) );
  NAND2X2 \mul/mult_6/U1236  ( .A(sig_B[9]), .B(sig_B[10]), .Y(
        \mul/mult_6/n666 ) );
  OAI21X1 \mul/mult_6/U1224  ( .A0(\mul/mult_6/n660 ), .A1(\mul/mult_6/n666 ), 
        .B0(\mul/mult_6/n661 ), .Y(\mul/mult_6/n659 ) );
  NOR2X2 \mul/mult_6/U1160  ( .A(\mul/mult_6/n620 ), .B(\mul/mult_6/n615 ), 
        .Y(\mul/mult_6/n613 ) );
  NOR2X2 \mul/mult_6/U1181  ( .A(\mul/mult_6/n635 ), .B(\mul/mult_6/n630 ), 
        .Y(\mul/mult_6/n628 ) );
  NOR2BX1 \mul/mult_6/U1069  ( .AN(\mul/mult_6/n1439 ), .B(\mul/mult_6/n1447 ), 
        .Y(\mul/mult_6/n531 ) );
  NOR2X2 \mul/mult_6/U1124  ( .A(\mul/mult_6/n596 ), .B(\mul/mult_6/n591 ), 
        .Y(\mul/mult_6/n589 ) );
  AOI21X1 \mul/mult_6/U1115  ( .A0(\mul/mult_6/n590 ), .A1(n592), .B0(
        \mul/mult_6/n585 ), .Y(\mul/mult_6/n583 ) );
  NAND2X2 \mul/mult_6/U1221  ( .A(\mul/mult_6/n670 ), .B(\mul/mult_6/n658 ), 
        .Y(\mul/mult_6/n652 ) );
  NOR2X2 \mul/mult_6/U1112  ( .A(\mul/mult_6/n599 ), .B(\mul/mult_6/n582 ), 
        .Y(\mul/mult_6/n580 ) );
  OAI21X1 \mul/mult_6/U572  ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1100 ), .Y(\mul/mult_6/n1074 ) );
  OAI21X1 \mul/mult_6/U745  ( .A0(n678), .A1(\mul/mult_6/n38 ), .B0(n531), .Y(
        \mul/mult_6/n1180 ) );
  OAI21X1 \mul/mult_6/U575  ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n58 ), 
        .B0(n535), .Y(\mul/mult_6/n1075 ) );
  OAI21XL \mul/mult_6/U984  ( .A0(n546), .A1(\mul/mult_6/n8 ), .B0(
        \mul/mult_6/n1359 ), .Y(\mul/mult_6/n1333 ) );
  OAI21X1 \mul/mult_6/U579  ( .A0(n678), .A1(\mul/mult_6/n58 ), .B0(n536), .Y(
        \mul/mult_6/n1076 ) );
  OAI21X1 \mul/mult_6/U655  ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1152 ), .Y(\mul/mult_6/n1126 ) );
  OAI21X1 \mul/mult_6/U569  ( .A0(n546), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1099 ), .Y(\mul/mult_6/n1073 ) );
  OAI21X1 \mul/mult_6/U652  ( .A0(n546), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1151 ), .Y(\mul/mult_6/n1125 ) );
  OAI21X1 \mul/mult_6/U658  ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n48 ), 
        .B0(n527), .Y(\mul/mult_6/n1127 ) );
  OAI21X1 \mul/mult_6/U662  ( .A0(n678), .A1(\mul/mult_6/n48 ), .B0(n530), .Y(
        \mul/mult_6/n1128 ) );
  XOR2X1 \mul/mult_6/U827  ( .A(\mul/mult_6/n1232 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n892 ) );
  XOR2X1 \mul/mult_6/U823  ( .A(\mul/mult_6/n1231 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n891 ) );
  XOR2X1 \mul/mult_6/U906  ( .A(\mul/mult_6/n1283 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n918 ) );
  XOR2X1 \mul/mult_6/U910  ( .A(\mul/mult_6/n1284 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n919 ) );
  XOR2XL \mul/mult_6/U986  ( .A(\mul/mult_6/n1334 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n944 ) );
  XOR2X1 \mul/mult_6/U661  ( .A(\mul/mult_6/n1128 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n838 ) );
  XOR2X1 \mul/mult_6/U654  ( .A(\mul/mult_6/n1126 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n836 ) );
  XOR2X1 \mul/mult_6/U820  ( .A(\mul/mult_6/n1230 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n890 ) );
  OAI21X1 \mul/mult_6/U1248  ( .A0(\mul/mult_6/n677 ), .A1(\mul/mult_6/n675 ), 
        .B0(\mul/mult_6/n676 ), .Y(\mul/mult_6/n674 ) );
  XOR2X1 \mul/mult_6/U734  ( .A(\mul/mult_6/n1177 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n862 ) );
  XOR2X1 \mul/mult_6/U657  ( .A(\mul/mult_6/n1127 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n837 ) );
  ADDFX1 \expadd/add_0_root_sub_0_root_sub_8/U4  ( .A(\expadd/N5 ), .B(
        exp_B[5]), .CI(\expadd/add_0_root_sub_0_root_sub_8/n5 ), .CO(
        \expadd/add_0_root_sub_0_root_sub_8/n4 ), .S(exp_P[5]) );
  XOR2X1 \mul/mult_6/U744  ( .A(\mul/mult_6/n1180 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n865 ) );
  XOR2X1 \mul/mult_6/U737  ( .A(\mul/mult_6/n1178 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n863 ) );
  XOR2X1 \mul/mult_6/U740  ( .A(\mul/mult_6/n1179 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n864 ) );
  XOR2X1 \mul/mult_6/U817  ( .A(\mul/mult_6/n1229 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n889 ) );
  XOR2X1 \mul/mult_6/U651  ( .A(\mul/mult_6/n1125 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n835 ) );
  CLKNAND2X2 \mul/mult_6/U180  ( .A(\mul/mult_6/n946 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n175 ) );
  XOR2X1 \mul/mult_6/U731  ( .A(\mul/mult_6/n1176 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n861 ) );
  ADDFX1 \expadd/add_0_root_sub_0_root_sub_8/U3  ( .A(\expadd/N6 ), .B(
        exp_B[6]), .CI(\expadd/add_0_root_sub_0_root_sub_8/n4 ), .CO(
        \expadd/add_0_root_sub_0_root_sub_8/n3 ), .S(exp_P[6]) );
  ADDHX1 \mul/mult_6/U295  ( .A(sig_A[14]), .B(\mul/mult_6/n838 ), .CO(
        \mul/mult_6/n461 ), .S(\mul/mult_6/n462 ) );
  AOI21X1 \mul/mult_6/U1131  ( .A0(\mul/mult_6/n598 ), .A1(\mul/mult_6/n713 ), 
        .B0(\mul/mult_6/n595 ), .Y(\mul/mult_6/n593 ) );
  OAI21X1 \mul/mult_6/U670  ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1182 ), .Y(\mul/mult_6/n1156 ) );
  XOR2X1 \mul/mult_6/U648  ( .A(\mul/mult_6/n1124 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n834 ) );
  XOR2X1 \mul/mult_6/U897  ( .A(\mul/mult_6/n1280 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n915 ) );
  AOI21X1 \mul/mult_6/U1123  ( .A0(\mul/mult_6/n598 ), .A1(\mul/mult_6/n589 ), 
        .B0(\mul/mult_6/n590 ), .Y(\mul/mult_6/n588 ) );
  XOR2X1 \mul/mult_6/U1174  ( .A(\mul/mult_6/n632 ), .B(\mul/mult_6/n559 ), 
        .Y(\mul/mult_6/n1398 ) );
  OAI21X1 \mul/mult_6/U750  ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n28 ), 
        .B0(n684), .Y(\mul/mult_6/n1207 ) );
  OAI21X1 \mul/mult_6/U809  ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1252 ), .Y(\mul/mult_6/n1226 ) );
  OAI21X1 \mul/mult_6/U465  ( .A0(n542), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1040 ), .Y(\mul/mult_6/n1014 ) );
  XOR2X1 \mul/mult_6/U1138  ( .A(\mul/mult_6/n605 ), .B(\mul/mult_6/n555 ), 
        .Y(\mul/mult_6/n1394 ) );
  OAI21X1 \mul/mult_6/U435  ( .A0(n591), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1030 ), .Y(\mul/mult_6/n1004 ) );
  OAI21X1 \mul/mult_6/U542  ( .A0(n572), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1090 ), .Y(\mul/mult_6/n1064 ) );
  OAI21X1 \mul/mult_6/U667  ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n38 ), 
        .B0(n686), .Y(\mul/mult_6/n1155 ) );
  OAI21X1 \mul/mult_6/U601  ( .A0(n591), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1134 ), .Y(\mul/mult_6/n1108 ) );
  OAI21X1 \mul/mult_6/U524  ( .A0(n569), .A1(\mul/mult_6/n58 ), .B0(
        \mul/mult_6/n1084 ), .Y(\mul/mult_6/n1058 ) );
  OAI21X1 \mul/mult_6/U726  ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1200 ), .Y(\mul/mult_6/n1174 ) );
  OAI21X1 \mul/mult_6/U613  ( .A0(n570), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1138 ), .Y(\mul/mult_6/n1112 ) );
  OAI21X1 \mul/mult_6/U607  ( .A0(n569), .A1(\mul/mult_6/n48 ), .B0(
        \mul/mult_6/n1136 ), .Y(\mul/mult_6/n1110 ) );
  XOR2X1 \mul/mult_6/U1215  ( .A(\mul/mult_6/n662 ), .B(\mul/mult_6/n563 ), 
        .Y(\mul/mult_6/n1402 ) );
  OAI21X1 \mul/mult_6/U643  ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1148 ), .Y(\mul/mult_6/n1122 ) );
  XOR2X1 \mul/mult_6/U1156  ( .A(\mul/mult_6/n617 ), .B(\mul/mult_6/n557 ), 
        .Y(\mul/mult_6/n1396 ) );
  XOR2X1 \mul/mult_6/U811  ( .A(\mul/mult_6/n1227 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n887 ) );
  XOR2X1 \mul/mult_6/U796  ( .A(\mul/mult_6/n1222 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n882 ) );
  ADDFX1 \mul/mult_6/U198  ( .A(n672), .B(\mul/mult_6/n217 ), .CI(n652), .CO(
        \mul/mult_6/n211 ), .S(\mul/mult_6/n212 ) );
  XOR2X1 \mul/mult_6/U639  ( .A(\mul/mult_6/n1121 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n831 ) );
  XOR2X1 \mul/mult_6/U722  ( .A(\mul/mult_6/n1173 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n858 ) );
  XOR2X1 \mul/mult_6/U950  ( .A(\mul/mult_6/n1322 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n932 ) );
  XOR2X1 \mul/mult_6/U808  ( .A(\mul/mult_6/n1226 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n886 ) );
  XOR2X1 \mul/mult_6/U805  ( .A(\mul/mult_6/n1225 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n885 ) );
  XOR2X1 \mul/mult_6/U956  ( .A(\mul/mult_6/n1324 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n934 ) );
  ADDFX1 \mul/mult_6/U217  ( .A(n675), .B(\mul/mult_6/n266 ), .CI(n642), .CO(
        \mul/mult_6/n257 ), .S(\mul/mult_6/n258 ) );
  XOR2X1 \mul/mult_6/U891  ( .A(\mul/mult_6/n1278 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n913 ) );
  XOR2X1 \mul/mult_6/U790  ( .A(\mul/mult_6/n1220 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n880 ) );
  XOR2X1 \mul/mult_6/U645  ( .A(\mul/mult_6/n1123 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n833 ) );
  XOR2X1 \mul/mult_6/U944  ( .A(\mul/mult_6/n1320 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n930 ) );
  XOR2X1 \mul/mult_6/U867  ( .A(\mul/mult_6/n1270 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n905 ) );
  XOR2X1 \mul/mult_6/U725  ( .A(\mul/mult_6/n1174 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n859 ) );
  XOR2X1 \mul/mult_6/U642  ( .A(\mul/mult_6/n1122 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n832 ) );
  XOR2X1 \mul/mult_6/U873  ( .A(\mul/mult_6/n1272 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n907 ) );
  XOR2X1 \mul/mult_6/U630  ( .A(\mul/mult_6/n1118 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n828 ) );
  XOR2X1 \mul/mult_6/U728  ( .A(\mul/mult_6/n1175 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n860 ) );
  XOR2X1 \mul/mult_6/U802  ( .A(\mul/mult_6/n1224 ), .B(sig_A[8]), .Y(
        \mul/mult_6/n884 ) );
  OAI21X1 \mul/mult_6/U512  ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1080 ), .Y(\mul/mult_6/n1054 ) );
  OAI21X1 \mul/mult_6/U533  ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1087 ), .Y(\mul/mult_6/n1061 ) );
  OAI21X1 \mul/mult_6/U438  ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1031 ), .Y(\mul/mult_6/n1005 ) );
  OAI21X1 \mul/mult_6/U456  ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1037 ), .Y(\mul/mult_6/n1011 ) );
  ADDFX1 \mul/mult_6/U302  ( .A(\mul/mult_6/n481 ), .B(\mul/mult_6/n938 ), 
        .CI(\mul/mult_6/n914 ), .CO(\mul/mult_6/n478 ), .S(\mul/mult_6/n479 )
         );
  ADDFX1 \mul/mult_6/U249  ( .A(sig_B[1]), .B(n605), .CI(\mul/mult_6/n353 ), 
        .CO(\mul/mult_6/n342 ), .S(\mul/mult_6/n343 ) );
  OAI21X1 \mul/mult_6/U595  ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1132 ), .Y(\mul/mult_6/n1106 ) );
  ADDFX1 \mul/mult_6/U213  ( .A(sig_B[10]), .B(n675), .CI(\mul/mult_6/n768 ), 
        .CO(\mul/mult_6/n248 ), .S(\mul/mult_6/n249 ) );
  OAI21X1 \mul/mult_6/U545  ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1091 ), .Y(\mul/mult_6/n1065 ) );
  OAI21X1 \mul/mult_6/U840  ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1287 ), .Y(\mul/mult_6/n1261 ) );
  OAI21X1 \mul/mult_6/U521  ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1083 ), .Y(\mul/mult_6/n1057 ) );
  OAI21X1 \mul/mult_6/U444  ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1033 ), .Y(\mul/mult_6/n1007 ) );
  OAI21X1 \mul/mult_6/U515  ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1081 ), .Y(\mul/mult_6/n1055 ) );
  OAI21X1 \mul/mult_6/U610  ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1137 ), .Y(\mul/mult_6/n1111 ) );
  OAI21X1 \mul/mult_6/U757  ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1235 ), .Y(\mul/mult_6/n1209 ) );
  OAI21X1 \mul/mult_6/U462  ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n68 ), 
        .B0(\mul/mult_6/n1039 ), .Y(\mul/mult_6/n1013 ) );
  OAI21X1 \mul/mult_6/U508  ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n58 ), 
        .B0(\mul/mult_6/n1079 ), .Y(\mul/mult_6/n1053 ) );
  OAI21X1 \mul/mult_6/U598  ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n48 ), 
        .B0(\mul/mult_6/n1133 ), .Y(\mul/mult_6/n1107 ) );
  XOR2X1 \mul/mult_6/U947  ( .A(\mul/mult_6/n1321 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n931 ) );
  XOR2X1 \mul/mult_6/U953  ( .A(\mul/mult_6/n1323 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n933 ) );
  XOR2X1 \mul/mult_6/U876  ( .A(\mul/mult_6/n1273 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n908 ) );
  MXI2X1 \align/sra_11/U583  ( .A(\align/sra_11/n475 ), .B(\align/sra_11/n476 ), .S0(n719), .Y(\align/sra_11/n473 ) );
  MXI2X1 \align/sra_11/U579  ( .A(\align/sra_11/n468 ), .B(\align/sra_11/n469 ), .S0(n719), .Y(\align/sra_11/n466 ) );
  MXI2X1 \align/sra_11/U724  ( .A(\align/sra_11/n736 ), .B(\align/sra_11/n595 ), .S0(n719), .Y(\align/sra_11/n731 ) );
  MXI2X1 \align/sra_11/U713  ( .A(\align/sra_11/n729 ), .B(\align/sra_11/n591 ), .S0(n719), .Y(\align/sra_11/n728 ) );
  ADDFX2 \mul/mult_6/U158  ( .A(\mul/mult_6/n420 ), .B(\mul/mult_6/n427 ), 
        .CI(\mul/mult_6/n158 ), .CO(\mul/mult_6/n157 ), .S(sig_P[17]) );
  ADDFX2 \mul/mult_6/U157  ( .A(\mul/mult_6/n410 ), .B(\mul/mult_6/n419 ), 
        .CI(\mul/mult_6/n157 ), .CO(\mul/mult_6/n156 ), .S(sig_P[18]) );
  MXI2XL \align/sra_11/U641  ( .A(\align/sra_11/n586 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n585 ) );
  MXI2XL \align/sra_11/U639  ( .A(\align/sra_11/n582 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n581 ) );
  MXI2XL \align/sra_11/U654  ( .A(\align/sra_11/n615 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n614 ) );
  MXI2XL \align/sra_11/U434  ( .A(\align/sra_11/n556 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n555 ) );
  MXI2XL \align/sra_11/U647  ( .A(\align/sra_11/n598 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n597 ) );
  MXI2XL \align/sra_11/U631  ( .A(\align/sra_11/n566 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n565 ) );
  MXI2XL \align/sra_11/U658  ( .A(\align/sra_11/n621 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n620 ) );
  MXI2XL \align/sra_11/U676  ( .A(\align/sra_11/n655 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n654 ) );
  MXI2XL \align/sra_11/U626  ( .A(\align/sra_11/n558 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n557 ) );
  MXI2XL \align/sra_11/U645  ( .A(\align/sra_11/n594 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n593 ) );
  MXI2XL \align/sra_11/U629  ( .A(\align/sra_11/n562 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n561 ) );
  MXI2XL \align/sra_11/U662  ( .A(\align/sra_11/n627 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n626 ) );
  MXI2XL \align/sra_11/U672  ( .A(\align/sra_11/n649 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n648 ) );
  MXI2XL \align/sra_11/U424  ( .A(\align/sra_11/n603 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n602 ) );
  MXI2XL \align/sra_11/U643  ( .A(\align/sra_11/n590 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n589 ) );
  MXI2XL \align/sra_11/U650  ( .A(\align/sra_11/n609 ), .B(\two_en[1] ), .S0(
        n717), .Y(\align/sra_11/n608 ) );
  MXI2XL \align/sra_11/U668  ( .A(\align/sra_11/n643 ), .B(\two_en[1] ), .S0(
        n515), .Y(\align/sra_11/n642 ) );
  MXI2X1 \align/sra_11/U632  ( .A(n722), .B(\align/sra_11/n569 ), .S0(n510), 
        .Y(\align/N56 ) );
  MXI2X1 \align/sra_10/U331  ( .A(sel_P[22]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n277 ) );
  MXI2XL \align/sra_10/U353  ( .A(sig_P[0]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n255 ) );
  MXI2X2 \align/sra_10/U304  ( .A(n707), .B(n706), .S0(n509), .Y(
        \align/sra_10/n304 ) );
  MXI2X2 \align/sra_10/U305  ( .A(sel_P[48]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n303 ) );
  MXI2X1 \align/sra_10/U248  ( .A(\align/sra_10/n202 ), .B(\align/sra_10/n204 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n152 ) );
  MXI2X1 \align/sra_10/U58  ( .A(\align/sra_10/n92 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n42 ) );
  MXI2X1 \align/sra_10/U98  ( .A(\align/sra_10/n52 ), .B(\align/sra_10/n84 ), 
        .S0(n717), .Y(\align/sra_10/n2 ) );
  MXI2X1 \align/sra_10/U57  ( .A(\align/sra_10/n93 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n43 ) );
  MXI2X1 \align/sra_10/U52  ( .A(\align/sra_10/n98 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n48 ) );
  MXI2X1 \align/sra_10/U53  ( .A(\align/sra_10/n97 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n47 ) );
  MXI2X1 \align/sra_10/U96  ( .A(\align/sra_10/n54 ), .B(\align/sra_10/n86 ), 
        .S0(n717), .Y(\align/sra_10/n4 ) );
  MXI2X1 \align/sra_10/U54  ( .A(\align/sra_10/n96 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n46 ) );
  MXI2X1 \align/sra_10/U97  ( .A(\align/sra_10/n53 ), .B(\align/sra_10/n85 ), 
        .S0(n717), .Y(\align/sra_10/n3 ) );
  MXI2X1 \align/sra_10/U56  ( .A(\align/sra_10/n94 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n44 ) );
  MXI2X1 \align/sra_10/U55  ( .A(\align/sra_10/n95 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n45 ) );
  MXI2X1 \align/sra_10/U51  ( .A(\align/sra_10/n99 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n49 ) );
  MX2X1 \align/sra_10/U49  ( .A(\align/sra_10/n1 ), .B(\align/sra_10/n17 ), 
        .S0(n719), .Y(\align/N4 ) );
  MX2X1 \align/sra_10/U16  ( .A(\align/sra_10/n34 ), .B(\align/sra_10/n50 ), 
        .S0(n718), .Y(\align/N37 ) );
  MX2X1 \align/sra_10/U15  ( .A(\align/sra_10/n35 ), .B(n706), .S0(n718), .Y(
        \align/N38 ) );
  MX2X1 \align/sra_10/U19  ( .A(\align/sra_10/n31 ), .B(\align/sra_10/n47 ), 
        .S0(n718), .Y(\align/N34 ) );
  MX2X1 \align/sra_10/U17  ( .A(\align/sra_10/n33 ), .B(\align/sra_10/n49 ), 
        .S0(n718), .Y(\align/N36 ) );
  MX2X1 \align/sra_10/U24  ( .A(\align/sra_10/n26 ), .B(\align/sra_10/n42 ), 
        .S0(n718), .Y(\align/N29 ) );
  MX2X1 \align/sra_10/U20  ( .A(\align/sra_10/n30 ), .B(\align/sra_10/n46 ), 
        .S0(n718), .Y(\align/N33 ) );
  MX2X1 \align/sra_10/U18  ( .A(\align/sra_10/n32 ), .B(\align/sra_10/n48 ), 
        .S0(n718), .Y(\align/N35 ) );
  MX2X1 \align/sra_10/U23  ( .A(\align/sra_10/n27 ), .B(\align/sra_10/n43 ), 
        .S0(n718), .Y(\align/N30 ) );
  MX2X1 \align/sra_10/U21  ( .A(\align/sra_10/n29 ), .B(\align/sra_10/n45 ), 
        .S0(n718), .Y(\align/N32 ) );
  MX2X1 \align/sra_10/U22  ( .A(\align/sra_10/n28 ), .B(\align/sra_10/n44 ), 
        .S0(n718), .Y(\align/N31 ) );
  NAND2X2 \sigadd/add_9/U243  ( .A(ali_P[15]), .B(ali_C[15]), .Y(
        \sigadd/add_9/n188 ) );
  NAND2X2 \sigadd/add_9/U117  ( .A(ali_P[33]), .B(ali_C[33]), .Y(
        \sigadd/add_9/n116 ) );
  NAND2X2 \sigadd/add_9/U229  ( .A(ali_P[17]), .B(ali_C[17]), .Y(
        \sigadd/add_9/n180 ) );
  NAND2X2 \sigadd/add_9/U103  ( .A(ali_P[35]), .B(ali_C[35]), .Y(
        \sigadd/add_9/n108 ) );
  NAND2X2 \sigadd/add_9/U223  ( .A(ali_P[18]), .B(ali_C[18]), .Y(
        \sigadd/add_9/n177 ) );
  NAND2X2 \sigadd/add_9/U131  ( .A(ali_P[31]), .B(ali_C[31]), .Y(
        \sigadd/add_9/n124 ) );
  NAND2X2 \sigadd/add_9/U187  ( .A(ali_P[23]), .B(ali_C[23]), .Y(
        \sigadd/add_9/n156 ) );
  NAND2X2 \sigadd/add_9/U201  ( .A(ali_P[21]), .B(ali_C[21]), .Y(
        \sigadd/add_9/n164 ) );
  NAND2X2 \sigadd/add_9/U215  ( .A(ali_P[19]), .B(ali_C[19]), .Y(
        \sigadd/add_9/n172 ) );
  NAND2X2 \sigadd/add_9/U145  ( .A(ali_P[29]), .B(ali_C[29]), .Y(
        \sigadd/add_9/n132 ) );
  NAND2X2 \sigadd/add_9/U159  ( .A(ali_P[27]), .B(ali_C[27]), .Y(
        \sigadd/add_9/n140 ) );
  NAND2X2 \sigadd/add_9/U173  ( .A(ali_P[25]), .B(ali_C[25]), .Y(
        \sigadd/add_9/n148 ) );
  CLKNAND2X2 \sigadd/add_9/U343  ( .A(n561), .B(\sigadd/add_9/n246 ), .Y(
        \sigadd/add_9/n50 ) );
  NAND2XL \sigadd/add_9/U338  ( .A(\sigadd/add_9/n295 ), .B(
        \sigadd/add_9/n244 ), .Y(\sigadd/add_9/n49 ) );
  MXI2XL \normal/srl_15/U235  ( .A(\normal/srl_15/n208 ), .B(
        \normal/srl_15/n210 ), .S0(n715), .Y(\normal/srl_15/n158 ) );
  MXI2XL \normal/sll_15/U190  ( .A(\normal/sll_15/n233 ), .B(
        \normal/sll_15/n231 ), .S0(n514), .Y(\normal/sll_15/n186 ) );
  MXI2XL \normal/srl_15/U234  ( .A(\normal/srl_15/n209 ), .B(
        \normal/srl_15/n211 ), .S0(n715), .Y(\normal/srl_15/n159 ) );
  MXI2XL \normal/sll_15/U188  ( .A(\normal/sll_15/n235 ), .B(
        \normal/sll_15/n233 ), .S0(n514), .Y(\normal/sll_15/n188 ) );
  MXI2XL \normal/srl_15/U233  ( .A(\normal/srl_15/n210 ), .B(
        \normal/srl_15/n212 ), .S0(n715), .Y(\normal/srl_15/n160 ) );
  MXI2XL \normal/sll_15/U191  ( .A(\normal/sll_15/n232 ), .B(
        \normal/sll_15/n230 ), .S0(n514), .Y(\normal/sll_15/n185 ) );
  MXI2X1 \normal/sll_15/U49  ( .A(\normal/sll_15/n92 ), .B(\normal/sll_15/n88 ), .S0(n704), .Y(\normal/sll_15/n45 ) );
  MXI2X1 \normal/sll_15/U51  ( .A(\normal/sll_15/n90 ), .B(\normal/sll_15/n86 ), .S0(n704), .Y(\normal/sll_15/n43 ) );
  MXI2X1 \normal/sll_15/U72  ( .A(\normal/sll_15/n69 ), .B(\normal/sll_15/n65 ), .S0(n704), .Y(\normal/sll_15/n22 ) );
  MXI2X1 \normal/sll_15/U50  ( .A(\normal/sll_15/n91 ), .B(\normal/sll_15/n87 ), .S0(n704), .Y(\normal/sll_15/n44 ) );
  MXI2X1 \normal/sll_15/U52  ( .A(\normal/sll_15/n89 ), .B(\normal/sll_15/n85 ), .S0(n704), .Y(\normal/sll_15/n42 ) );
  NOR2X2 \ctrl/add_1_root_add_16_2/U33  ( .A(n525), .B(
        \ctrl/add_1_root_add_16_2/n48 ), .Y(\ctrl/add_1_root_add_16_2/n30 ) );
  NAND2X2 \round/r298/U26  ( .A(norm_out[22]), .B(norm_out[23]), .Y(
        \round/r298/n21 ) );
  NAND2X2 \round/r298/U104  ( .A(norm_out[10]), .B(norm_out[11]), .Y(
        \round/r298/n87 ) );
  NAND2X2 \round/r298/U79  ( .A(norm_out[15]), .B(norm_out[14]), .Y(
        \round/r298/n66 ) );
  NAND2X2 \round/r298/U127  ( .A(norm_out[7]), .B(norm_out[6]), .Y(
        \round/r298/n106 ) );
  NAND2X2 \round/r298/U51  ( .A(norm_out[18]), .B(norm_out[19]), .Y(
        \round/r298/n42 ) );
  XOR2X1 \round/r298/U60  ( .A(\round/r298/n57 ), .B(\round/r298/n56 ), .Y(
        \round/N22 ) );
  XOR2X1 \round/r298/U15  ( .A(\round/r298/n17 ), .B(\round/r298/n16 ), .Y(
        \round/N29 ) );
  XOR2X1 \round/r298/U35  ( .A(\round/r298/n36 ), .B(\round/r298/n35 ), .Y(
        \round/N26 ) );
  XOR2X1 \round/r298/U47  ( .A(\round/r298/n45 ), .B(\round/r298/n44 ), .Y(
        \round/N24 ) );
  XOR2X1 \round/r298/U88  ( .A(\round/r298/n81 ), .B(\round/r298/n80 ), .Y(
        \round/N18 ) );
  XOR2X1 \round/r298/U54  ( .A(\round/r298/n50 ), .B(\round/r298/n49 ), .Y(
        \round/N23 ) );
  NAND2X2 \ctrl/sub_0_root_add_0_root_sub_16/U32  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[3] ), .B(n709), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n26 ) );
  XOR2X1 \ctrl/sub_0_root_add_0_root_sub_16/U41  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/n6 ), .B(
        \ctrl/sub_0_root_add_0_root_sub_16/n35 ), .Y(\ctrl/N28 ) );
  NOR2X4 \ctrl/sub_0_root_add_0_root_sub_16/U17  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[5] ), .B(n713), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n8 ) );
  XOR2X1 \ctrl/sub_0_root_add_0_root_sub_16/U27  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/n4 ), .B(
        \ctrl/sub_0_root_add_0_root_sub_16/n27 ), .Y(\ctrl/N30 ) );
  NOR2X2 \mul/mult_6/U1136  ( .A(sig_B[19]), .B(sig_B[20]), .Y(
        \mul/mult_6/n596 ) );
  NOR2X2 \mul/mult_6/U1172  ( .A(sig_B[15]), .B(sig_B[16]), .Y(
        \mul/mult_6/n620 ) );
  NOR2X2 \mul/mult_6/U1258  ( .A(\mul/mult_6/n686 ), .B(\mul/mult_6/n683 ), 
        .Y(\mul/mult_6/n681 ) );
  NOR2X2 \mul/mult_6/U1241  ( .A(\mul/mult_6/n675 ), .B(\mul/mult_6/n672 ), 
        .Y(\mul/mult_6/n670 ) );
  NOR2X2 \mul/mult_6/U1142  ( .A(\mul/mult_6/n608 ), .B(\mul/mult_6/n603 ), 
        .Y(\mul/mult_6/n601 ) );
  AO21XL \mul/mult_6/U344  ( .A0(n696), .A1(sig_B[22]), .B0(n695), .Y(
        \mul/mult_6/n520 ) );
  OAI21X1 \mul/mult_6/U828  ( .A0(n678), .A1(\mul/mult_6/n28 ), .B0(n532), .Y(
        \mul/mult_6/n1232 ) );
  OAI21X1 \mul/mult_6/U824  ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n28 ), 
        .B0(n529), .Y(\mul/mult_6/n1231 ) );
  OAI21X1 \mul/mult_6/U738  ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n38 ), 
        .B0(\mul/mult_6/n1204 ), .Y(\mul/mult_6/n1178 ) );
  OAI21X1 \mul/mult_6/U741  ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n38 ), 
        .B0(n528), .Y(\mul/mult_6/n1179 ) );
  OAI21X1 \mul/mult_6/U818  ( .A0(n546), .A1(\mul/mult_6/n28 ), .B0(
        \mul/mult_6/n1255 ), .Y(\mul/mult_6/n1229 ) );
  OAI21X1 \mul/mult_6/U735  ( .A0(n546), .A1(\mul/mult_6/n38 ), .B0(
        \mul/mult_6/n1203 ), .Y(\mul/mult_6/n1177 ) );
  OAI21X1 \mul/mult_6/U821  ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n28 ), 
        .B0(\mul/mult_6/n1256 ), .Y(\mul/mult_6/n1230 ) );
  XOR2X1 \mul/mult_6/U993  ( .A(\mul/mult_6/n1336 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n946 ) );
  XOR2X1 \mul/mult_6/U1264  ( .A(\mul/mult_6/n688 ), .B(\mul/mult_6/n568 ), 
        .Y(\mul/mult_6/n1407 ) );
  ADDHX1 \mul/mult_6/U301  ( .A(sig_A[11]), .B(\mul/mult_6/n865 ), .CO(
        \mul/mult_6/n476 ), .S(\mul/mult_6/n477 ) );
  ADDHX1 \mul/mult_6/U307  ( .A(sig_A[8]), .B(\mul/mult_6/n892 ), .CO(
        \mul/mult_6/n488 ), .S(\mul/mult_6/n489 ) );
  AOI21X1 \mul/mult_6/U1111  ( .A0(\mul/mult_6/n622 ), .A1(\mul/mult_6/n580 ), 
        .B0(\mul/mult_6/n581 ), .Y(\mul/mult_6/n579 ) );
  XOR2X1 \mul/mult_6/U1122  ( .A(\mul/mult_6/n593 ), .B(\mul/mult_6/n553 ), 
        .Y(\mul/mult_6/n1392 ) );
  XOR2X1 \mul/mult_6/U1110  ( .A(\mul/mult_6/n588 ), .B(\mul/mult_6/n552 ), 
        .Y(\mul/mult_6/n1391 ) );
  XOR2X1 \mul/mult_6/U1103  ( .A(\mul/mult_6/n579 ), .B(sig_B[22]), .Y(
        \mul/mult_6/n1390 ) );
  XOR2X1 \mul/mult_6/U968  ( .A(\mul/mult_6/n1328 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n938 ) );
  XOR2X1 \mul/mult_6/U888  ( .A(\mul/mult_6/n1277 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n912 ) );
  XOR2X1 \mul/mult_6/U965  ( .A(\mul/mult_6/n1327 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n937 ) );
  XOR2X1 \mul/mult_6/U962  ( .A(\mul/mult_6/n1326 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n936 ) );
  XOR2X1 \mul/mult_6/U882  ( .A(\mul/mult_6/n1275 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n910 ) );
  ADDFX1 \mul/mult_6/U268  ( .A(\mul/mult_6/n397 ), .B(\mul/mult_6/n830 ), 
        .CI(\mul/mult_6/n806 ), .CO(\mul/mult_6/n394 ), .S(\mul/mult_6/n395 )
         );
  XOR2X1 \mul/mult_6/U959  ( .A(\mul/mult_6/n1325 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n935 ) );
  ADDFX1 \mul/mult_6/U272  ( .A(\mul/mult_6/n407 ), .B(\mul/mult_6/n807 ), 
        .CI(\mul/mult_6/n414 ), .CO(\mul/mult_6/n404 ), .S(\mul/mult_6/n405 )
         );
  ADDFX2 \mul/mult_6/U159  ( .A(\mul/mult_6/n428 ), .B(\mul/mult_6/n435 ), 
        .CI(\mul/mult_6/n159 ), .CO(\mul/mult_6/n158 ), .S(sig_P[16]) );
  INVX2 \align/sra_11/U360  ( .A(\align/sra_11/n560 ), .Y(\align/sra_11/n757 )
         );
  MX2X1 \align/sra_11/U727  ( .A(\two_en[1] ), .B(\align/sra_11/n753 ), .S0(
        n510), .Y(\align/N54 ) );
  ADDFHX2 \mul/mult_6/U147  ( .A(\mul/mult_6/n302 ), .B(\mul/mult_6/n312 ), 
        .CI(\mul/mult_6/n147 ), .CO(\mul/mult_6/n146 ), .S(sig_P[28]) );
  ADDFHX2 \mul/mult_6/U145  ( .A(\mul/mult_6/n281 ), .B(\mul/mult_6/n290 ), 
        .CI(\mul/mult_6/n145 ), .CO(\mul/mult_6/n144 ), .S(sig_P[30]) );
  ADDFHX2 \mul/mult_6/U139  ( .A(\mul/mult_6/n235 ), .B(\mul/mult_6/n229 ), 
        .CI(\mul/mult_6/n139 ), .CO(\mul/mult_6/n138 ), .S(sig_P[36]) );
  ADDFHX2 \mul/mult_6/U136  ( .A(\mul/mult_6/n215 ), .B(\mul/mult_6/n210 ), 
        .CI(\mul/mult_6/n136 ), .CO(\mul/mult_6/n135 ), .S(sig_P[39]) );
  ADDFHX2 \mul/mult_6/U135  ( .A(\mul/mult_6/n209 ), .B(\mul/mult_6/n204 ), 
        .CI(\mul/mult_6/n135 ), .CO(\mul/mult_6/n134 ), .S(sig_P[40]) );
  ADDFHX2 \mul/mult_6/U134  ( .A(\mul/mult_6/n203 ), .B(\mul/mult_6/n199 ), 
        .CI(\mul/mult_6/n134 ), .CO(\mul/mult_6/n133 ), .S(sig_P[41]) );
  ADDFHX2 \mul/mult_6/U133  ( .A(\mul/mult_6/n198 ), .B(\mul/mult_6/n195 ), 
        .CI(\mul/mult_6/n133 ), .CO(\mul/mult_6/n132 ), .S(sig_P[42]) );
  MXI2X1 \align/sra_10/U316  ( .A(sel_P[37]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n292 ) );
  MXI2X1 \align/sra_10/U329  ( .A(sel_P[24]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n279 ) );
  MXI2X1 \align/sra_10/U312  ( .A(sel_P[41]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n296 ) );
  MXI2X1 \align/sra_10/U319  ( .A(sel_P[34]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n289 ) );
  MXI2X1 \align/sra_10/U318  ( .A(sel_P[35]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n290 ) );
  MXI2X1 \align/sra_10/U323  ( .A(sel_P[30]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n285 ) );
  MXI2X1 \align/sra_10/U314  ( .A(sel_P[39]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n294 ) );
  MXI2X1 \align/sra_10/U324  ( .A(sel_P[29]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n284 ) );
  MXI2X1 \align/sra_10/U308  ( .A(sel_P[45]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n300 ) );
  MXI2X1 \align/sra_10/U307  ( .A(sel_P[46]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n301 ) );
  MXI2X1 \align/sra_10/U326  ( .A(sel_P[27]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n282 ) );
  MXI2X1 \align/sra_10/U317  ( .A(sel_P[36]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n291 ) );
  MXI2X1 \align/sra_10/U309  ( .A(sel_P[44]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n299 ) );
  MXI2X1 \align/sra_10/U313  ( .A(sel_P[40]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n295 ) );
  MXI2X1 \align/sra_10/U311  ( .A(sel_P[42]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n297 ) );
  MXI2X1 \align/sra_10/U327  ( .A(sel_P[26]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n281 ) );
  MXI2X1 \align/sra_10/U320  ( .A(sel_P[33]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n288 ) );
  MXI2X1 \align/sra_10/U322  ( .A(sel_P[31]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n286 ) );
  MXI2X1 \align/sra_10/U321  ( .A(sel_P[32]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n287 ) );
  MXI2X1 \align/sra_10/U315  ( .A(sel_P[38]), .B(n707), .S0(n509), .Y(
        \align/sra_10/n293 ) );
  NAND2XL \sigadd/add_9/U5  ( .A(n706), .B(\two_en[1] ), .Y(\sigadd/add_9/n52 ) );
  MXI2X1 \align/sra_10/U306  ( .A(sel_P[47]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n302 ) );
  MXI2X1 \align/sra_10/U310  ( .A(sel_P[43]), .B(n706), .S0(n509), .Y(
        \align/sra_10/n298 ) );
  MXI2X2 \align/sra_10/U250  ( .A(\align/sra_10/n304 ), .B(n508), .S0(n507), 
        .Y(\align/sra_10/n250 ) );
  MXI2X1 \align/sra_10/U208  ( .A(\align/sra_10/n242 ), .B(\align/sra_10/n244 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n192 ) );
  MXI2X1 \align/sra_10/U213  ( .A(\align/sra_10/n237 ), .B(\align/sra_10/n239 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n187 ) );
  MXI2X1 \align/sra_10/U210  ( .A(\align/sra_10/n240 ), .B(\align/sra_10/n242 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n190 ) );
  MXI2X1 \align/sra_10/U216  ( .A(\align/sra_10/n234 ), .B(\align/sra_10/n236 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n184 ) );
  MXI2X1 \align/sra_10/U209  ( .A(\align/sra_10/n241 ), .B(\align/sra_10/n243 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n191 ) );
  MXI2X1 \align/sra_10/U212  ( .A(\align/sra_10/n238 ), .B(\align/sra_10/n240 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n188 ) );
  MXI2X1 \align/sra_10/U220  ( .A(\align/sra_10/n230 ), .B(\align/sra_10/n232 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n180 ) );
  MXI2X1 \align/sra_10/U226  ( .A(\align/sra_10/n224 ), .B(\align/sra_10/n226 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n174 ) );
  MXI2X1 \align/sra_10/U211  ( .A(\align/sra_10/n239 ), .B(\align/sra_10/n241 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n189 ) );
  MXI2X1 \align/sra_10/U225  ( .A(\align/sra_10/n225 ), .B(\align/sra_10/n227 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n175 ) );
  MXI2X1 \align/sra_10/U205  ( .A(\align/sra_10/n245 ), .B(\align/sra_10/n247 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n195 ) );
  MXI2X1 \align/sra_10/U204  ( .A(\align/sra_10/n246 ), .B(\align/sra_10/n248 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n196 ) );
  MXI2X1 \align/sra_10/U206  ( .A(\align/sra_10/n244 ), .B(\align/sra_10/n246 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n194 ) );
  MXI2X1 \align/sra_10/U218  ( .A(\align/sra_10/n232 ), .B(\align/sra_10/n234 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n182 ) );
  MXI2X1 \align/sra_10/U249  ( .A(\align/sra_10/n201 ), .B(\align/sra_10/n203 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n151 ) );
  MXI2X1 \align/sra_10/U173  ( .A(\align/sra_10/n177 ), .B(\align/sra_10/n181 ), .S0(n505), .Y(\align/sra_10/n127 ) );
  MXI2X1 \align/sra_10/U180  ( .A(\align/sra_10/n170 ), .B(\align/sra_10/n174 ), .S0(n505), .Y(\align/sra_10/n120 ) );
  MXI2X1 \align/sra_10/U177  ( .A(\align/sra_10/n173 ), .B(\align/sra_10/n177 ), .S0(n505), .Y(\align/sra_10/n123 ) );
  MXI2X1 \align/sra_10/U181  ( .A(\align/sra_10/n169 ), .B(\align/sra_10/n173 ), .S0(n505), .Y(\align/sra_10/n119 ) );
  MXI2X1 \align/sra_10/U199  ( .A(\align/sra_10/n151 ), .B(\align/sra_10/n155 ), .S0(n505), .Y(\align/sra_10/n101 ) );
  MXI2X1 \align/sra_10/U169  ( .A(\align/sra_10/n181 ), .B(\align/sra_10/n185 ), .S0(n511), .Y(\align/sra_10/n131 ) );
  MXI2X1 \align/sra_10/U179  ( .A(\align/sra_10/n171 ), .B(\align/sra_10/n175 ), .S0(n505), .Y(\align/sra_10/n121 ) );
  MXI2X1 \align/sra_10/U178  ( .A(\align/sra_10/n172 ), .B(\align/sra_10/n176 ), .S0(n505), .Y(\align/sra_10/n122 ) );
  MXI2X1 \align/sra_10/U168  ( .A(\align/sra_10/n182 ), .B(\align/sra_10/n186 ), .S0(n511), .Y(\align/sra_10/n132 ) );
  MXI2X1 \align/sra_10/U176  ( .A(\align/sra_10/n174 ), .B(\align/sra_10/n178 ), .S0(n505), .Y(\align/sra_10/n124 ) );
  MXI2X1 \align/sra_10/U175  ( .A(\align/sra_10/n175 ), .B(\align/sra_10/n179 ), .S0(n511), .Y(\align/sra_10/n125 ) );
  MXI2X1 \align/sra_10/U171  ( .A(\align/sra_10/n179 ), .B(\align/sra_10/n183 ), .S0(n511), .Y(\align/sra_10/n129 ) );
  MXI2X1 \align/sra_10/U110  ( .A(\align/sra_10/n140 ), .B(\align/sra_10/n148 ), .S0(n705), .Y(\align/sra_10/n90 ) );
  MXI2X1 \align/sra_10/U107  ( .A(\align/sra_10/n143 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n93 ) );
  MXI2X1 \align/sra_10/U102  ( .A(\align/sra_10/n148 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n98 ) );
  MXI2X1 \align/sra_10/U149  ( .A(\align/sra_10/n101 ), .B(\align/sra_10/n109 ), .S0(n506), .Y(\align/sra_10/n51 ) );
  MXI2X1 \align/sra_10/U103  ( .A(\align/sra_10/n147 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n97 ) );
  MXI2X1 \align/sra_10/U105  ( .A(\align/sra_10/n145 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n95 ) );
  MXI2X1 \align/sra_10/U101  ( .A(\align/sra_10/n149 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n99 ) );
  MXI2X1 \align/sra_10/U106  ( .A(\align/sra_10/n144 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n94 ) );
  MXI2X1 \align/sra_10/U104  ( .A(\align/sra_10/n146 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n96 ) );
  MXI2X1 \align/sra_10/U109  ( .A(\align/sra_10/n141 ), .B(\align/sra_10/n149 ), .S0(n705), .Y(\align/sra_10/n91 ) );
  MXI2X1 \align/sra_10/U108  ( .A(\align/sra_10/n142 ), .B(\align/sra_10/n150 ), .S0(n705), .Y(\align/sra_10/n92 ) );
  MXI2X1 \align/sra_10/U111  ( .A(\align/sra_10/n139 ), .B(\align/sra_10/n147 ), .S0(n705), .Y(\align/sra_10/n89 ) );
  MXI2X1 \align/sra_10/U112  ( .A(\align/sra_10/n138 ), .B(\align/sra_10/n146 ), .S0(n705), .Y(\align/sra_10/n88 ) );
  MXI2X1 \align/sra_10/U115  ( .A(\align/sra_10/n135 ), .B(\align/sra_10/n143 ), .S0(n705), .Y(\align/sra_10/n85 ) );
  MXI2X1 \align/sra_10/U113  ( .A(\align/sra_10/n137 ), .B(\align/sra_10/n145 ), .S0(n705), .Y(\align/sra_10/n87 ) );
  MXI2X1 \align/sra_10/U116  ( .A(\align/sra_10/n134 ), .B(\align/sra_10/n142 ), .S0(n705), .Y(\align/sra_10/n84 ) );
  MXI2X1 \align/sra_10/U100  ( .A(\align/sra_10/n150 ), .B(n706), .S0(n705), 
        .Y(\align/sra_10/n100 ) );
  MXI2X1 \align/sra_10/U114  ( .A(\align/sra_10/n136 ), .B(\align/sra_10/n144 ), .S0(n705), .Y(\align/sra_10/n86 ) );
  MXI2X1 \align/sra_10/U81  ( .A(\align/sra_10/n69 ), .B(n508), .S0(n717), .Y(
        \align/sra_10/n19 ) );
  MXI2X1 \align/sra_10/U65  ( .A(\align/sra_10/n85 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n35 ) );
  MXI2X1 \align/sra_10/U69  ( .A(\align/sra_10/n81 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n31 ) );
  MXI2X1 \align/sra_10/U74  ( .A(\align/sra_10/n76 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n26 ) );
  MXI2X1 \align/sra_10/U99  ( .A(\align/sra_10/n51 ), .B(\align/sra_10/n83 ), 
        .S0(n515), .Y(\align/sra_10/n1 ) );
  MXI2X1 \align/sra_10/U64  ( .A(\align/sra_10/n86 ), .B(n508), .S0(n717), .Y(
        \align/sra_10/n36 ) );
  MXI2X1 \align/sra_10/U79  ( .A(\align/sra_10/n71 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n21 ) );
  MXI2X1 \align/sra_10/U66  ( .A(\align/sra_10/n84 ), .B(n508), .S0(n717), .Y(
        \align/sra_10/n34 ) );
  MXI2X1 \align/sra_10/U75  ( .A(\align/sra_10/n75 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n25 ) );
  MXI2X1 \align/sra_10/U62  ( .A(\align/sra_10/n88 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n38 ) );
  MXI2X1 \align/sra_10/U72  ( .A(\align/sra_10/n78 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n28 ) );
  MXI2X1 \align/sra_10/U63  ( .A(\align/sra_10/n87 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n37 ) );
  MXI2X1 \align/sra_10/U70  ( .A(\align/sra_10/n80 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n30 ) );
  MXI2X1 \align/sra_10/U67  ( .A(\align/sra_10/n83 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n33 ) );
  MXI2X1 \align/sra_10/U68  ( .A(\align/sra_10/n82 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n32 ) );
  MXI2X1 \align/sra_10/U71  ( .A(\align/sra_10/n79 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n29 ) );
  MXI2X1 \align/sra_10/U78  ( .A(\align/sra_10/n72 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n22 ) );
  MXI2X1 \align/sra_10/U59  ( .A(\align/sra_10/n91 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n41 ) );
  MXI2X1 \align/sra_10/U60  ( .A(\align/sra_10/n90 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n40 ) );
  MXI2X1 \align/sra_10/U76  ( .A(\align/sra_10/n74 ), .B(n508), .S0(n717), .Y(
        \align/sra_10/n24 ) );
  MXI2X1 \align/sra_10/U77  ( .A(\align/sra_10/n73 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n23 ) );
  MXI2X1 \align/sra_10/U61  ( .A(\align/sra_10/n89 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n39 ) );
  MXI2X1 \align/sra_10/U80  ( .A(\align/sra_10/n70 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n20 ) );
  MXI2X1 \align/sra_10/U73  ( .A(\align/sra_10/n77 ), .B(n508), .S0(n515), .Y(
        \align/sra_10/n27 ) );
  MX2X1 \align/sra_10/U27  ( .A(\align/sra_10/n23 ), .B(\align/sra_10/n39 ), 
        .S0(n718), .Y(\align/N26 ) );
  MX2X1 \align/sra_10/U26  ( .A(\align/sra_10/n24 ), .B(\align/sra_10/n40 ), 
        .S0(n718), .Y(\align/N27 ) );
  MX2XL \align/sra_10/U3  ( .A(\align/sra_10/n47 ), .B(n706), .S0(n718), .Y(
        \align/N50 ) );
  MX2X1 \align/sra_10/U28  ( .A(\align/sra_10/n22 ), .B(\align/sra_10/n38 ), 
        .S0(n718), .Y(\align/N25 ) );
  MX2X1 \align/sra_10/U30  ( .A(\align/sra_10/n20 ), .B(\align/sra_10/n36 ), 
        .S0(n718), .Y(\align/N23 ) );
  MX2XL \align/sra_10/U1  ( .A(\align/sra_10/n49 ), .B(n706), .S0(n718), .Y(
        \align/N52 ) );
  MX2X1 \align/sra_10/U31  ( .A(\align/sra_10/n19 ), .B(\align/sra_10/n35 ), 
        .S0(n718), .Y(\align/N22 ) );
  MX2X1 \align/sra_10/U29  ( .A(\align/sra_10/n21 ), .B(\align/sra_10/n37 ), 
        .S0(n718), .Y(\align/N24 ) );
  MX2XL \align/sra_10/U4  ( .A(\align/sra_10/n46 ), .B(n706), .S0(n718), .Y(
        \align/N49 ) );
  MX2X1 \align/sra_10/U25  ( .A(\align/sra_10/n25 ), .B(\align/sra_10/n41 ), 
        .S0(n718), .Y(\align/N28 ) );
  MX2XL \align/sra_10/U2  ( .A(\align/sra_10/n48 ), .B(n706), .S0(n718), .Y(
        \align/N51 ) );
  NOR2X2 \sigadd/add_9/U18  ( .A(ali_P[47]), .B(ali_C[47]), .Y(
        \sigadd/add_9/n59 ) );
  NOR2X2 \sigadd/add_9/U46  ( .A(ali_P[43]), .B(ali_C[43]), .Y(
        \sigadd/add_9/n75 ) );
  NOR2X2 \sigadd/add_9/U74  ( .A(ali_P[39]), .B(ali_C[39]), .Y(
        \sigadd/add_9/n91 ) );
  NOR2X2 \sigadd/add_9/U102  ( .A(ali_P[35]), .B(ali_C[35]), .Y(
        \sigadd/add_9/n107 ) );
  NOR2X2 \sigadd/add_9/U32  ( .A(ali_P[45]), .B(ali_C[45]), .Y(
        \sigadd/add_9/n67 ) );
  NOR2X2 \sigadd/add_9/U88  ( .A(ali_P[37]), .B(ali_C[37]), .Y(
        \sigadd/add_9/n99 ) );
  NOR2X2 \sigadd/add_9/U60  ( .A(ali_P[41]), .B(ali_C[41]), .Y(
        \sigadd/add_9/n83 ) );
  OAI21X2 \sigadd/add_9/U337  ( .A0(\sigadd/add_9/n243 ), .A1(
        \sigadd/add_9/n246 ), .B0(\sigadd/add_9/n244 ), .Y(\sigadd/add_9/n242 ) );
  OAI21X4 \sigadd/add_9/U323  ( .A0(\sigadd/add_9/n237 ), .A1(
        \sigadd/add_9/n235 ), .B0(\sigadd/add_9/n236 ), .Y(\sigadd/add_9/n234 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U25  ( .A(n615), .B(\sigadd/sub_add_11_b0/n25 ), 
        .CO(\sigadd/sub_add_11_b0/n24 ), .S(\sigadd/N27 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U22  ( .A(n602), .B(\sigadd/sub_add_11_b0/n22 ), 
        .CO(\sigadd/sub_add_11_b0/n21 ), .S(\sigadd/N30 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U21  ( .A(n613), .B(\sigadd/sub_add_11_b0/n21 ), 
        .CO(\sigadd/sub_add_11_b0/n20 ), .S(\sigadd/N31 ) );
  MXI2XL \normal/sll_15/U189  ( .A(\normal/sll_15/n234 ), .B(
        \normal/sll_15/n232 ), .S0(n514), .Y(\normal/sll_15/n187 ) );
  MXI2X1 \normal/sll_15/U59  ( .A(\normal/sll_15/n82 ), .B(\normal/sll_15/n78 ), .S0(n704), .Y(\normal/sll_15/n35 ) );
  MXI2X1 \normal/sll_15/U48  ( .A(\normal/sll_15/n93 ), .B(\normal/sll_15/n89 ), .S0(n704), .Y(\normal/sll_15/n46 ) );
  MXI2X1 \normal/srl_15/U72  ( .A(\normal/srl_15/n71 ), .B(\normal/srl_15/n75 ), .S0(n704), .Y(\normal/srl_15/n23 ) );
  MXI2X1 \normal/sll_15/U53  ( .A(\normal/sll_15/n88 ), .B(\normal/sll_15/n84 ), .S0(n704), .Y(\normal/sll_15/n41 ) );
  MXI2X1 \normal/sll_15/U58  ( .A(\normal/sll_15/n83 ), .B(\normal/sll_15/n79 ), .S0(n704), .Y(\normal/sll_15/n36 ) );
  MXI2X1 \normal/sll_15/U71  ( .A(\normal/sll_15/n70 ), .B(\normal/sll_15/n66 ), .S0(\normal/n30 ), .Y(\normal/sll_15/n23 ) );
  MXI2X1 \normal/sll_15/U54  ( .A(\normal/sll_15/n87 ), .B(\normal/sll_15/n83 ), .S0(n704), .Y(\normal/sll_15/n40 ) );
  MXI2X1 \normal/sll_15/U24  ( .A(\normal/sll_15/n24 ), .B(\normal/sll_15/n23 ), .S0(n503), .Y(\normal/N71 ) );
  MXI2X1 \normal/srl_15/U24  ( .A(\normal/srl_15/n24 ), .B(\normal/srl_15/n25 ), .S0(n503), .Y(\normal/N25 ) );
  MXI2X1 \normal/sll_15/U1  ( .A(\normal/sll_15/n47 ), .B(\normal/sll_15/n46 ), 
        .S0(n503), .Y(\normal/N94 ) );
  MXI2X1 \normal/srl_15/U25  ( .A(\normal/srl_15/n23 ), .B(\normal/srl_15/n24 ), .S0(n503), .Y(\normal/N24 ) );
  MXI2X1 \normal/sll_15/U25  ( .A(\normal/sll_15/n23 ), .B(\normal/sll_15/n22 ), .S0(n503), .Y(\normal/N70 ) );
  NOR2X4 \round/r298/U78  ( .A(\round/r298/n66 ), .B(\round/r298/n76 ), .Y(
        \round/r298/n63 ) );
  NAND2X2 \round/r298/U12  ( .A(norm_out[25]), .B(norm_out[24]), .Y(
        \round/r298/n9 ) );
  NOR2X2 \round/r298/U50  ( .A(\round/r298/n52 ), .B(\round/r298/n42 ), .Y(
        \round/r298/n41 ) );
  NOR2X2 \round/r298/U7  ( .A(\round/r298/n9 ), .B(n556), .Y(\round/r298/n5 )
         );
  AOI21X1 \ctrl/add_1_root_add_16_2/U70  ( .A0(n702), .A1(n520), .B0(
        \ctrl/add_1_root_add_16_2/n60 ), .Y(\ctrl/add_1_root_add_16_2/n58 ) );
  AOI21X1 \ctrl/add_1_root_add_16_2/U44  ( .A0(n702), .A1(
        \ctrl/add_1_root_add_16_2/n39 ), .B0(\ctrl/add_1_root_add_16_2/n40 ), 
        .Y(\ctrl/add_1_root_add_16_2/n38 ) );
  OAI21X2 \ctrl/sub_0_root_add_0_root_sub_16/U42  ( .A0(
        \ctrl/sub_0_root_add_0_root_sub_16/n33 ), .A1(
        \ctrl/sub_0_root_add_0_root_sub_16/n35 ), .B0(
        \ctrl/sub_0_root_add_0_root_sub_16/n34 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n32 ) );
  NAND2X2 \ctrl/sub_0_root_add_0_root_sub_16/U26  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[4] ), .B(n708), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n23 ) );
  NOR2X2 \mul/mult_6/U1154  ( .A(sig_B[17]), .B(sig_B[18]), .Y(
        \mul/mult_6/n608 ) );
  NOR2X2 \mul/mult_6/U1235  ( .A(sig_B[9]), .B(sig_B[10]), .Y(
        \mul/mult_6/n665 ) );
  NOR2X2 \mul/mult_6/U1223  ( .A(\mul/mult_6/n665 ), .B(\mul/mult_6/n660 ), 
        .Y(\mul/mult_6/n658 ) );
  XNOR2XL \sub/sub_17/U10  ( .A(\expadd/add_0_root_sub_0_root_sub_8/n2 ), .B(
        exp_C[0]), .Y(\sub/N14 ) );
  XNOR2XL \sub/r301/U10  ( .A(exp_P[0]), .B(\sub/r301/n17 ), .Y(\sub/N5 ) );
  AO21XL \mul/mult_6/U427  ( .A0(n693), .A1(sig_B[22]), .B0(n692), .Y(
        \mul/mult_6/n524 ) );
  AO21XL \mul/mult_6/U676  ( .A0(n698), .A1(sig_B[22]), .B0(n685), .Y(
        \mul/mult_6/n536 ) );
  OAI21X1 \mul/mult_6/U1178  ( .A0(\mul/mult_6/n653 ), .A1(\mul/mult_6/n626 ), 
        .B0(\mul/mult_6/n627 ), .Y(\mul/mult_6/n625 ) );
  OAI21X1 \mul/mult_6/U901  ( .A0(n546), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1307 ), .Y(\mul/mult_6/n1281 ) );
  OAI21XL \mul/mult_6/U994  ( .A0(n678), .A1(\mul/mult_6/n8 ), .B0(n524), .Y(
        \mul/mult_6/n1336 ) );
  XOR2X1 \mul/mult_6/U900  ( .A(\mul/mult_6/n1281 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n916 ) );
  OAI21X1 \mul/mult_6/U898  ( .A0(n545), .A1(\mul/mult_6/n18 ), .B0(
        \mul/mult_6/n1306 ), .Y(\mul/mult_6/n1280 ) );
  XOR2X1 \mul/mult_6/U903  ( .A(\mul/mult_6/n1282 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n917 ) );
  AOI21X1 \mul/mult_6/U1167  ( .A0(\mul/mult_6/n622 ), .A1(\mul/mult_6/n717 ), 
        .B0(\mul/mult_6/n619 ), .Y(\mul/mult_6/n617 ) );
  AOI21X1 \mul/mult_6/U1149  ( .A0(\mul/mult_6/n610 ), .A1(\mul/mult_6/n715 ), 
        .B0(\mul/mult_6/n607 ), .Y(\mul/mult_6/n605 ) );
  AOI21X1 \mul/mult_6/U1188  ( .A0(\mul/mult_6/n637 ), .A1(\mul/mult_6/n719 ), 
        .B0(\mul/mult_6/n634 ), .Y(\mul/mult_6/n632 ) );
  OAI21X1 \mul/mult_6/U895  ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1305 ), .Y(\mul/mult_6/n1279 ) );
  CLKNAND2X2 \mul/mult_6/U177  ( .A(n640), .B(\mul/mult_6/n175 ), .Y(
        \mul/mult_6/n125 ) );
  XOR2XL \mul/mult_6/U586  ( .A(\mul/mult_6/n1104 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n814 ) );
  OAI21X1 \mul/mult_6/U892  ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1304 ), .Y(\mul/mult_6/n1278 ) );
  XOR2X1 \mul/mult_6/U894  ( .A(\mul/mult_6/n1279 ), .B(sig_A[5]), .Y(
        \mul/mult_6/n914 ) );
  XOR2X1 \mul/mult_6/U971  ( .A(\mul/mult_6/n1329 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n939 ) );
  XOR2XL \mul/mult_6/U583  ( .A(\mul/mult_6/n1103 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n813 ) );
  XOR2XL \mul/mult_6/U590  ( .A(\mul/mult_6/n1105 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n815 ) );
  XOR2XL \mul/mult_6/U428  ( .A(\mul/mult_6/n1002 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n762 ) );
  ADDHX1 \selc/r299/U9  ( .A(\selc/r299/n9 ), .B(\selc/r299/A[41] ), .CO(
        \selc/r299/n8 ), .S(\selc/N154 ) );
  ADDHX1 \selc/r299/U8  ( .A(\selc/r299/n8 ), .B(\selc/r299/A[42] ), .CO(
        \selc/r299/n7 ), .S(\selc/N155 ) );
  ADDHX1 \selc/r299/U7  ( .A(\selc/r299/n7 ), .B(\selc/r299/A[43] ), .CO(
        \selc/r299/n6 ), .S(\selc/N156 ) );
  ADDHX1 \selc/r299/U6  ( .A(\selc/r299/n6 ), .B(\selc/r299/A[44] ), .CO(
        \selc/r299/n5 ), .S(\selc/N157 ) );
  ADDHX2 \selc/r299/U5  ( .A(\selc/r299/n5 ), .B(\selc/r299/A[45] ), .CO(
        \selc/r299/n4 ), .S(\selc/N158 ) );
  ADDHX2 \selc/r299/U4  ( .A(\selc/r299/n4 ), .B(\selc/r299/A[46] ), .CO(
        \selc/r299/n3 ), .S(\selc/N159 ) );
  XOR2X4 \selc/r299/U1  ( .A(\selc/r299/n1 ), .B(\mul/mult_6/n126 ), .Y(
        \selc/N162 ) );
  MXI2X1 \align/sra_10/U265  ( .A(\align/sra_10/n289 ), .B(\align/sra_10/n290 ), .S0(n507), .Y(\align/sra_10/n235 ) );
  MXI2X1 \align/sra_10/U215  ( .A(\align/sra_10/n235 ), .B(\align/sra_10/n237 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n185 ) );
  MXI2X1 \align/sra_10/U207  ( .A(\align/sra_10/n243 ), .B(\align/sra_10/n245 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n193 ) );
  MXI2X1 \align/sra_10/U214  ( .A(\align/sra_10/n236 ), .B(\align/sra_10/n238 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n186 ) );
  MXI2X1 \align/sra_10/U221  ( .A(\align/sra_10/n229 ), .B(\align/sra_10/n231 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n179 ) );
  MXI2X1 \align/sra_10/U222  ( .A(\align/sra_10/n228 ), .B(\align/sra_10/n230 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n178 ) );
  MXI2X1 \align/sra_10/U223  ( .A(\align/sra_10/n227 ), .B(\align/sra_10/n229 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n177 ) );
  MXI2X1 \align/sra_10/U202  ( .A(\align/sra_10/n248 ), .B(\align/sra_10/n250 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n198 ) );
  MXI2X1 \align/sra_10/U227  ( .A(\align/sra_10/n223 ), .B(\align/sra_10/n225 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n173 ) );
  MXI2X1 \align/sra_10/U219  ( .A(\align/sra_10/n231 ), .B(\align/sra_10/n233 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n181 ) );
  MXI2X1 \align/sra_10/U203  ( .A(\align/sra_10/n247 ), .B(\align/sra_10/n249 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n197 ) );
  MXI2X1 \align/sra_10/U172  ( .A(\align/sra_10/n178 ), .B(\align/sra_10/n182 ), .S0(n511), .Y(\align/sra_10/n128 ) );
  MXI2X1 \align/sra_10/U163  ( .A(\align/sra_10/n187 ), .B(\align/sra_10/n191 ), .S0(n511), .Y(\align/sra_10/n137 ) );
  MXI2X1 \align/sra_10/U170  ( .A(\align/sra_10/n180 ), .B(\align/sra_10/n184 ), .S0(n511), .Y(\align/sra_10/n130 ) );
  MXI2X1 \align/sra_10/U164  ( .A(\align/sra_10/n186 ), .B(\align/sra_10/n190 ), .S0(n511), .Y(\align/sra_10/n136 ) );
  MX2X1 \align/sra_10/U34  ( .A(\align/sra_10/n16 ), .B(\align/sra_10/n32 ), 
        .S0(n718), .Y(\align/N19 ) );
  MX2XL \align/sra_10/U5  ( .A(\align/sra_10/n45 ), .B(n706), .S0(n718), .Y(
        \align/N48 ) );
  MX2X1 \align/sra_10/U40  ( .A(\align/sra_10/n10 ), .B(\align/sra_10/n26 ), 
        .S0(n718), .Y(\align/N13 ) );
  MX2X1 \align/sra_10/U35  ( .A(\align/sra_10/n15 ), .B(\align/sra_10/n31 ), 
        .S0(n718), .Y(\align/N18 ) );
  MX2XL \align/sra_10/U6  ( .A(\align/sra_10/n44 ), .B(n706), .S0(n718), .Y(
        \align/N47 ) );
  MX2X1 \align/sra_10/U38  ( .A(\align/sra_10/n12 ), .B(\align/sra_10/n28 ), 
        .S0(n718), .Y(\align/N15 ) );
  MX2X1 \align/sra_10/U39  ( .A(\align/sra_10/n11 ), .B(\align/sra_10/n27 ), 
        .S0(n718), .Y(\align/N14 ) );
  MX2X1 \align/sra_10/U36  ( .A(\align/sra_10/n14 ), .B(\align/sra_10/n30 ), 
        .S0(n718), .Y(\align/N17 ) );
  MX2X1 \align/sra_10/U37  ( .A(\align/sra_10/n13 ), .B(\align/sra_10/n29 ), 
        .S0(n718), .Y(\align/N16 ) );
  MX2XL \align/sra_10/U8  ( .A(\align/sra_10/n42 ), .B(n706), .S0(n718), .Y(
        \align/N45 ) );
  MX2X1 \align/sra_10/U32  ( .A(\align/sra_10/n18 ), .B(\align/sra_10/n34 ), 
        .S0(n718), .Y(\align/N21 ) );
  MX2X1 \align/sra_10/U42  ( .A(\align/sra_10/n8 ), .B(\align/sra_10/n24 ), 
        .S0(n718), .Y(\align/N11 ) );
  MX2X1 \align/sra_10/U43  ( .A(\align/sra_10/n7 ), .B(\align/sra_10/n23 ), 
        .S0(n718), .Y(\align/N10 ) );
  MX2X1 \align/sra_10/U41  ( .A(\align/sra_10/n9 ), .B(\align/sra_10/n25 ), 
        .S0(n718), .Y(\align/N12 ) );
  MX2XL \align/sra_10/U7  ( .A(\align/sra_10/n43 ), .B(n706), .S0(n718), .Y(
        \align/N46 ) );
  MX2X1 \align/sra_10/U33  ( .A(\align/sra_10/n17 ), .B(\align/sra_10/n33 ), 
        .S0(n718), .Y(\align/N20 ) );
  NOR2X2 \sigadd/add_9/U158  ( .A(ali_P[27]), .B(ali_C[27]), .Y(
        \sigadd/add_9/n139 ) );
  NOR2X2 \sigadd/add_9/U186  ( .A(ali_P[23]), .B(ali_C[23]), .Y(
        \sigadd/add_9/n155 ) );
  NOR2X2 \sigadd/add_9/U172  ( .A(ali_P[25]), .B(ali_C[25]), .Y(
        \sigadd/add_9/n147 ) );
  NOR2X2 \sigadd/add_9/U116  ( .A(ali_P[33]), .B(ali_C[33]), .Y(
        \sigadd/add_9/n115 ) );
  NOR2X2 \sigadd/add_9/U130  ( .A(ali_P[31]), .B(ali_C[31]), .Y(
        \sigadd/add_9/n123 ) );
  NOR2X2 \sigadd/add_9/U144  ( .A(ali_P[29]), .B(ali_C[29]), .Y(
        \sigadd/add_9/n131 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U26  ( .A(n604), .B(\sigadd/sub_add_11_b0/n26 ), 
        .CO(\sigadd/sub_add_11_b0/n25 ), .S(\sigadd/N26 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U10  ( .A(n581), .B(\sigadd/sub_add_11_b0/n10 ), 
        .CO(\sigadd/sub_add_11_b0/n9 ), .S(\sigadd/N42 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U9  ( .A(n587), .B(\sigadd/sub_add_11_b0/n9 ), 
        .CO(\sigadd/sub_add_11_b0/n8 ), .S(\sigadd/N43 ) );
  ADDHX2 \sigadd/sub_add_11_b0/U8  ( .A(n580), .B(\sigadd/sub_add_11_b0/n8 ), 
        .CO(\sigadd/sub_add_11_b0/n7 ), .S(\sigadd/N44 ) );
  MXI2XL \normal/srl_15/U232  ( .A(\normal/srl_15/n211 ), .B(
        \normal/srl_15/n213 ), .S0(n715), .Y(\normal/srl_15/n161 ) );
  NOR2X1 \round/r298/U84  ( .A(\round/r298/n76 ), .B(\round/r298/n73 ), .Y(
        \round/r298/n70 ) );
  NAND2XL \round/r298/U22  ( .A(\round/r298/n1 ), .B(\round/r298/n18 ), .Y(
        \round/r298/n17 ) );
  AOI21X1 \ctrl/add_1_root_add_16_2/U12  ( .A0(n702), .A1(
        \ctrl/add_1_root_add_16_2/n16 ), .B0(\ctrl/add_1_root_add_16_2/n17 ), 
        .Y(\ctrl/add_1_root_add_16_2/n15 ) );
  AOI21X1 \ctrl/add_1_root_add_16_2/U4  ( .A0(n702), .A1(n526), .B0(n585), .Y(
        \ctrl/add_1_root_add_16_2/n8 ) );
  CLKXOR2X2 \mul/mult_6/U1059  ( .A(sig_A[19]), .B(sig_A[20]), .Y(
        \mul/mult_6/n1453 ) );
  AOI21X1 \mul/mult_6/U505  ( .A0(\mul/mult_6/n60 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n54 ), .Y(\mul/mult_6/n1078 ) );
  AOI21X1 \mul/mult_6/U422  ( .A0(\mul/mult_6/n70 ), .A1(sig_B[22]), .B0(
        \mul/mult_6/n64 ), .Y(\mul/mult_6/n1026 ) );
  AOI21X1 \mul/mult_6/U1257  ( .A0(\mul/mult_6/n681 ), .A1(\mul/mult_6/n690 ), 
        .B0(\mul/mult_6/n682 ), .Y(\mul/mult_6/n680 ) );
  ADDFXL \sub/r301/U8  ( .A(n659), .B(n1028), .CI(exp_P[1]), .CO(\sub/r301/n7 ), .S(\sub/N6 ) );
  ADDFXL \sub/sub_17/U8  ( .A(n660), .B(exp_C[1]), .CI(n1045), .CO(
        \sub/sub_17/n7 ), .S(\sub/N15 ) );
  OAI21X1 \mul/mult_6/U907  ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n18 ), 
        .B0(n564), .Y(\mul/mult_6/n1283 ) );
  OAI21X1 \mul/mult_6/U904  ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n18 ), 
        .B0(\mul/mult_6/n1308 ), .Y(\mul/mult_6/n1282 ) );
  AOI21X1 \mul/mult_6/U1230  ( .A0(\mul/mult_6/n667 ), .A1(\mul/mult_6/n723 ), 
        .B0(\mul/mult_6/n664 ), .Y(\mul/mult_6/n662 ) );
  AOI21X1 \mul/mult_6/U1208  ( .A0(\mul/mult_6/n651 ), .A1(\mul/mult_6/n721 ), 
        .B0(\mul/mult_6/n648 ), .Y(\mul/mult_6/n646 ) );
  CLKXOR2X2 \expadd/add_0_root_sub_0_root_sub_8/U1  ( .A(
        \expadd/add_0_root_sub_0_root_sub_8/n3 ), .B(
        \expadd/add_0_root_sub_0_root_sub_8/n1 ), .Y(exp_P[7]) );
  OAI21X1 \mul/mult_6/U975  ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1356 ), .Y(\mul/mult_6/n1330 ) );
  XOR2XL \mul/mult_6/U440  ( .A(\mul/mult_6/n1006 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n766 ) );
  XOR2X1 \mul/mult_6/U974  ( .A(\mul/mult_6/n1330 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n940 ) );
  XOR2X1 \mul/mult_6/U977  ( .A(\mul/mult_6/n1331 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n941 ) );
  XOR2XL \mul/mult_6/U915  ( .A(\mul/mult_6/n1311 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n921 ) );
  XOR2XL \mul/mult_6/U683  ( .A(\mul/mult_6/n1160 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n845 ) );
  XOR2XL \mul/mult_6/U695  ( .A(\mul/mult_6/n1164 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n849 ) );
  XOR2XL \sub/r301/U2  ( .A(exp_P[7]), .B(n1027), .Y(\sub/r301/n1 ) );
  XOR2XL \mul/mult_6/U449  ( .A(\mul/mult_6/n1009 ), .B(sig_A[20]), .Y(
        \mul/mult_6/n769 ) );
  XOR2XL \mul/mult_6/U677  ( .A(\mul/mult_6/n1158 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n843 ) );
  XOR2XL \mul/mult_6/U680  ( .A(\mul/mult_6/n1159 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n844 ) );
  XOR2XL \mul/mult_6/U673  ( .A(\mul/mult_6/n1157 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n842 ) );
  NOR2X1 \align/sra_11/U363  ( .A(sub_out[6]), .B(sub_out[7]), .Y(
        \align/sra_11/n465 ) );
  ADDFX2 \mul/mult_6/U165  ( .A(\mul/mult_6/n470 ), .B(\mul/mult_6/n474 ), 
        .CI(\mul/mult_6/n165 ), .CO(\mul/mult_6/n164 ), .S(sig_P[10]) );
  ADDFX2 \mul/mult_6/U164  ( .A(\mul/mult_6/n465 ), .B(\mul/mult_6/n469 ), 
        .CI(\mul/mult_6/n164 ), .CO(\mul/mult_6/n163 ), .S(sig_P[11]) );
  ADDFX2 \mul/mult_6/U156  ( .A(\mul/mult_6/n400 ), .B(\mul/mult_6/n409 ), 
        .CI(\mul/mult_6/n156 ), .CO(\mul/mult_6/n155 ), .S(sig_P[19]) );
  ADDFX2 \mul/mult_6/U130  ( .A(\mul/mult_6/n187 ), .B(\mul/mult_6/n184 ), 
        .CI(\mul/mult_6/n130 ), .CO(\mul/mult_6/n129 ), .S(sig_P[45]) );
  ADDFX2 \mul/mult_6/U129  ( .A(\mul/mult_6/n181 ), .B(\mul/mult_6/n183 ), 
        .CI(\mul/mult_6/n129 ), .CO(\mul/mult_6/n128 ), .S(sig_P[46]) );
  MXI2X1 \align/sra_10/U268  ( .A(\align/sra_10/n286 ), .B(\align/sra_10/n287 ), .S0(n507), .Y(\align/sra_10/n232 ) );
  MXI2X1 \align/sra_10/U272  ( .A(\align/sra_10/n282 ), .B(\align/sra_10/n283 ), .S0(n507), .Y(\align/sra_10/n228 ) );
  MXI2X1 \align/sra_10/U267  ( .A(\align/sra_10/n287 ), .B(\align/sra_10/n288 ), .S0(n507), .Y(\align/sra_10/n233 ) );
  MXI2X1 \align/sra_10/U263  ( .A(\align/sra_10/n291 ), .B(\align/sra_10/n292 ), .S0(n507), .Y(\align/sra_10/n237 ) );
  MXI2X1 \align/sra_10/U257  ( .A(\align/sra_10/n297 ), .B(\align/sra_10/n298 ), .S0(n507), .Y(\align/sra_10/n243 ) );
  MXI2X1 \align/sra_10/U275  ( .A(\align/sra_10/n279 ), .B(\align/sra_10/n280 ), .S0(n507), .Y(\align/sra_10/n225 ) );
  MXI2X1 \align/sra_10/U253  ( .A(\align/sra_10/n301 ), .B(\align/sra_10/n302 ), .S0(n507), .Y(\align/sra_10/n247 ) );
  MXI2X1 \align/sra_10/U269  ( .A(\align/sra_10/n285 ), .B(\align/sra_10/n286 ), .S0(n507), .Y(\align/sra_10/n231 ) );
  MXI2X1 \align/sra_10/U251  ( .A(\align/sra_10/n303 ), .B(\align/sra_10/n304 ), .S0(n507), .Y(\align/sra_10/n249 ) );
  MXI2X1 \align/sra_10/U255  ( .A(\align/sra_10/n299 ), .B(\align/sra_10/n300 ), .S0(n507), .Y(\align/sra_10/n245 ) );
  MXI2X1 \align/sra_10/U274  ( .A(\align/sra_10/n280 ), .B(\align/sra_10/n281 ), .S0(n507), .Y(\align/sra_10/n226 ) );
  MXI2X1 \align/sra_10/U259  ( .A(\align/sra_10/n295 ), .B(\align/sra_10/n296 ), .S0(n507), .Y(\align/sra_10/n241 ) );
  MXI2X1 \align/sra_10/U270  ( .A(\align/sra_10/n284 ), .B(\align/sra_10/n285 ), .S0(n507), .Y(\align/sra_10/n230 ) );
  MXI2X1 \align/sra_10/U277  ( .A(\align/sra_10/n277 ), .B(\align/sra_10/n278 ), .S0(n507), .Y(\align/sra_10/n223 ) );
  MXI2X1 \align/sra_10/U271  ( .A(\align/sra_10/n283 ), .B(\align/sra_10/n284 ), .S0(n507), .Y(\align/sra_10/n229 ) );
  MXI2X1 \align/sra_10/U261  ( .A(\align/sra_10/n293 ), .B(\align/sra_10/n294 ), .S0(n507), .Y(\align/sra_10/n239 ) );
  MXI2X1 \align/sra_10/U273  ( .A(\align/sra_10/n281 ), .B(\align/sra_10/n282 ), .S0(n507), .Y(\align/sra_10/n227 ) );
  MXI2X1 \align/sra_10/U229  ( .A(\align/sra_10/n221 ), .B(\align/sra_10/n223 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n171 ) );
  MXI2X1 \align/sra_10/U217  ( .A(\align/sra_10/n233 ), .B(\align/sra_10/n235 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n183 ) );
  MXI2X1 \align/sra_10/U224  ( .A(\align/sra_10/n226 ), .B(\align/sra_10/n228 ), .S0(\align/sra_11/SH[1] ), .Y(\align/sra_10/n176 ) );
  MXI2X1 \align/sra_10/U83  ( .A(\align/sra_10/n67 ), .B(\align/sra_10/n99 ), 
        .S0(n717), .Y(\align/sra_10/n17 ) );
  MX2XL \align/sra_10/U11  ( .A(\align/sra_10/n39 ), .B(n706), .S0(n718), .Y(
        \align/N42 ) );
  MX2XL \align/sra_10/U12  ( .A(\align/sra_10/n38 ), .B(n706), .S0(n718), .Y(
        \align/N41 ) );
  MX2XL \align/sra_10/U10  ( .A(\align/sra_10/n40 ), .B(n706), .S0(n718), .Y(
        \align/N43 ) );
  MX2XL \align/sra_10/U9  ( .A(\align/sra_10/n41 ), .B(n706), .S0(n718), .Y(
        \align/N44 ) );
  MX2XL \align/sra_10/U13  ( .A(\align/sra_10/n37 ), .B(n706), .S0(n718), .Y(
        \align/N40 ) );
  MX2XL \align/sra_10/U14  ( .A(\align/sra_10/n36 ), .B(n706), .S0(n718), .Y(
        \align/N39 ) );
  NOR2X2 \sigadd/add_9/U214  ( .A(ali_P[19]), .B(ali_C[19]), .Y(
        \sigadd/add_9/n171 ) );
  NOR2X2 \sigadd/add_9/U242  ( .A(ali_P[15]), .B(ali_C[15]), .Y(
        \sigadd/add_9/n187 ) );
  NOR2X2 \sigadd/add_9/U228  ( .A(ali_P[17]), .B(ali_C[17]), .Y(
        \sigadd/add_9/n179 ) );
  NOR2X2 \sigadd/add_9/U256  ( .A(ali_P[13]), .B(ali_C[13]), .Y(
        \sigadd/add_9/n195 ) );
  NOR2X2 \sigadd/add_9/U270  ( .A(ali_P[11]), .B(ali_C[11]), .Y(
        \sigadd/add_9/n203 ) );
  NOR2X2 \sigadd/add_9/U200  ( .A(ali_P[21]), .B(ali_C[21]), .Y(
        \sigadd/add_9/n163 ) );
  AOI21X4 \sigadd/add_9/U287  ( .A0(\sigadd/add_9/n218 ), .A1(n550), .B0(
        \sigadd/add_9/n215 ), .Y(\sigadd/add_9/n213 ) );
  OAI21X6 \sigadd/add_9/U253  ( .A0(\sigadd/add_9/n197 ), .A1(
        \sigadd/add_9/n195 ), .B0(\sigadd/add_9/n196 ), .Y(\sigadd/add_9/n194 ) );
  OAI21X6 \sigadd/add_9/U239  ( .A0(\sigadd/add_9/n189 ), .A1(
        \sigadd/add_9/n187 ), .B0(\sigadd/add_9/n188 ), .Y(\sigadd/add_9/n186 ) );
  AOI21X6 \sigadd/add_9/U231  ( .A0(\sigadd/add_9/n186 ), .A1(n579), .B0(
        \sigadd/add_9/n183 ), .Y(\sigadd/add_9/n181 ) );
  OAI21X6 \sigadd/add_9/U225  ( .A0(\sigadd/add_9/n181 ), .A1(
        \sigadd/add_9/n179 ), .B0(\sigadd/add_9/n180 ), .Y(\sigadd/add_9/n178 ) );
  AOI21X6 \sigadd/add_9/U217  ( .A0(\sigadd/add_9/n178 ), .A1(n578), .B0(
        \sigadd/add_9/n175 ), .Y(\sigadd/add_9/n173 ) );
  OAI21X6 \sigadd/add_9/U211  ( .A0(\sigadd/add_9/n173 ), .A1(
        \sigadd/add_9/n171 ), .B0(\sigadd/add_9/n172 ), .Y(\sigadd/add_9/n170 ) );
  OAI21X6 \sigadd/add_9/U197  ( .A0(\sigadd/add_9/n165 ), .A1(
        \sigadd/add_9/n163 ), .B0(\sigadd/add_9/n164 ), .Y(\sigadd/add_9/n162 ) );
  OAI21X6 \sigadd/add_9/U183  ( .A0(\sigadd/add_9/n157 ), .A1(
        \sigadd/add_9/n155 ), .B0(\sigadd/add_9/n156 ), .Y(\sigadd/add_9/n154 ) );
  OAI21X6 \sigadd/add_9/U169  ( .A0(\sigadd/add_9/n149 ), .A1(
        \sigadd/add_9/n147 ), .B0(\sigadd/add_9/n148 ), .Y(\sigadd/add_9/n146 ) );
  OAI21X6 \sigadd/add_9/U155  ( .A0(\sigadd/add_9/n141 ), .A1(
        \sigadd/add_9/n139 ), .B0(\sigadd/add_9/n140 ), .Y(\sigadd/add_9/n138 ) );
  OAI21X6 \sigadd/add_9/U141  ( .A0(\sigadd/add_9/n133 ), .A1(
        \sigadd/add_9/n131 ), .B0(\sigadd/add_9/n132 ), .Y(\sigadd/add_9/n130 ) );
  OAI21X6 \sigadd/add_9/U127  ( .A0(\sigadd/add_9/n125 ), .A1(
        \sigadd/add_9/n123 ), .B0(\sigadd/add_9/n124 ), .Y(\sigadd/add_9/n122 ) );
  OAI21X6 \sigadd/add_9/U113  ( .A0(\sigadd/add_9/n117 ), .A1(
        \sigadd/add_9/n115 ), .B0(\sigadd/add_9/n116 ), .Y(\sigadd/add_9/n114 ) );
  OAI21X6 \sigadd/add_9/U99  ( .A0(\sigadd/add_9/n109 ), .A1(
        \sigadd/add_9/n107 ), .B0(\sigadd/add_9/n108 ), .Y(\sigadd/add_9/n106 ) );
  OAI21X6 \sigadd/add_9/U85  ( .A0(\sigadd/add_9/n101 ), .A1(
        \sigadd/add_9/n99 ), .B0(\sigadd/add_9/n100 ), .Y(\sigadd/add_9/n98 )
         );
  OAI21X6 \sigadd/add_9/U71  ( .A0(\sigadd/add_9/n93 ), .A1(\sigadd/add_9/n91 ), .B0(\sigadd/add_9/n92 ), .Y(\sigadd/add_9/n90 ) );
  AOI21X4 \sigadd/add_9/U35  ( .A0(\sigadd/add_9/n74 ), .A1(n619), .B0(
        \sigadd/add_9/n71 ), .Y(\sigadd/add_9/n69 ) );
  AOI21X4 \sigadd/add_9/U21  ( .A0(\sigadd/add_9/n66 ), .A1(n618), .B0(
        \sigadd/add_9/n63 ), .Y(\sigadd/add_9/n61 ) );
  OAI21X4 \sigadd/add_9/U15  ( .A0(\sigadd/add_9/n61 ), .A1(\sigadd/add_9/n59 ), .B0(\sigadd/add_9/n60 ), .Y(\sigadd/add_9/n58 ) );
  NAND2X1 \ctrl/add_1_root_add_16_2/U73  ( .A(n520), .B(
        \ctrl/add_1_root_add_16_2/n62 ), .Y(\ctrl/add_1_root_add_16_2/n6 ) );
  NOR2X2 \round/r298/U103  ( .A(\round/r298/n87 ), .B(\round/r298/n95 ), .Y(
        \round/r298/n86 ) );
  NAND2XL \round/r298/U44  ( .A(\round/r298/n1 ), .B(norm_out[20]), .Y(
        \round/r298/n36 ) );
  NOR2X2 \ctrl/sub_0_root_add_0_root_sub_16/U48  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[0] ), .B(n711), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n35 ) );
  XNOR2X1 \mul/mult_6/U1064  ( .A(sig_A[15]), .B(sig_A[16]), .Y(
        \mul/mult_6/n1446 ) );
  NOR2X2 \mul/mult_6/U1164  ( .A(sig_B[16]), .B(sig_B[17]), .Y(
        \mul/mult_6/n615 ) );
  CLKXOR2X2 \mul/mult_6/U1066  ( .A(sig_A[16]), .B(sig_A[17]), .Y(
        \mul/mult_6/n1454 ) );
  XNOR2X1 \mul/mult_6/U1050  ( .A(sig_A[21]), .B(sig_A[22]), .Y(
        \mul/mult_6/n1444 ) );
  XNOR2X1 \mul/mult_6/U1057  ( .A(sig_A[18]), .B(sig_A[19]), .Y(
        \mul/mult_6/n1445 ) );
  OAI21X1 \mul/mult_6/U1202  ( .A0(\mul/mult_6/n644 ), .A1(\mul/mult_6/n650 ), 
        .B0(\mul/mult_6/n645 ), .Y(\mul/mult_6/n643 ) );
  NOR2X2 \mul/mult_6/U1201  ( .A(\mul/mult_6/n649 ), .B(\mul/mult_6/n644 ), 
        .Y(\mul/mult_6/n640 ) );
  CLKXOR2X2 \mul/mult_6/U1080  ( .A(sig_A[10]), .B(sig_A[11]), .Y(
        \mul/mult_6/n1456 ) );
  XNOR2X2 \mul/mult_6/U1072  ( .A(sig_A[11]), .B(sig_A[12]), .Y(
        \mul/mult_6/n1439 ) );
  CLKXOR2X2 \mul/mult_6/U1073  ( .A(sig_A[13]), .B(sig_A[14]), .Y(
        \mul/mult_6/n1455 ) );
  CLKXOR2X2 \mul/mult_6/U1094  ( .A(sig_A[4]), .B(sig_A[5]), .Y(
        \mul/mult_6/n1458 ) );
  OAI21X1 \mul/mult_6/U1125  ( .A0(\mul/mult_6/n591 ), .A1(\mul/mult_6/n597 ), 
        .B0(\mul/mult_6/n592 ), .Y(\mul/mult_6/n590 ) );
  OAI21X1 \mul/mult_6/U1113  ( .A0(\mul/mult_6/n600 ), .A1(\mul/mult_6/n582 ), 
        .B0(\mul/mult_6/n583 ), .Y(\mul/mult_6/n581 ) );
  XOR2X1 \mul/mult_6/U980  ( .A(\mul/mult_6/n1332 ), .B(sig_A[2]), .Y(
        \mul/mult_6/n942 ) );
  OAI21XL \mul/mult_6/U474  ( .A0(n544), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1043 ), .Y(\mul/mult_6/n1017 ) );
  ADDFX1 \mul/mult_6/U183  ( .A(sig_B[22]), .B(n670), .CI(n540), .CO(
        \mul/mult_6/n180 ), .S(\mul/mult_6/n181 ) );
  XOR2XL \mul/mult_6/U615  ( .A(\mul/mult_6/n1113 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n823 ) );
  ADDFX2 \mul/mult_6/U166  ( .A(\mul/mult_6/n475 ), .B(\mul/mult_6/n478 ), 
        .CI(\mul/mult_6/n166 ), .CO(\mul/mult_6/n165 ), .S(sig_P[9]) );
  ADDFX2 \mul/mult_6/U155  ( .A(\mul/mult_6/n390 ), .B(\mul/mult_6/n399 ), 
        .CI(\mul/mult_6/n155 ), .CO(\mul/mult_6/n154 ), .S(sig_P[20]) );
  ADDFX2 \mul/mult_6/U149  ( .A(\mul/mult_6/n324 ), .B(\mul/mult_6/n334 ), 
        .CI(\mul/mult_6/n149 ), .CO(\mul/mult_6/n148 ), .S(sig_P[26]) );
  ADDFX2 \mul/mult_6/U146  ( .A(\mul/mult_6/n291 ), .B(\mul/mult_6/n301 ), 
        .CI(\mul/mult_6/n146 ), .CO(\mul/mult_6/n145 ), .S(sig_P[29]) );
  MXI2X1 \align/sra_10/U167  ( .A(\align/sra_10/n183 ), .B(\align/sra_10/n187 ), .S0(n511), .Y(\align/sra_10/n133 ) );
  NOR2X2 \normal/srl_15/U95  ( .A(\normal/srl_15/n148 ), .B(n513), .Y(
        \normal/srl_15/n98 ) );
  NOR2X2 \normal/srl_15/U96  ( .A(\normal/srl_15/n147 ), .B(n513), .Y(
        \normal/srl_15/n97 ) );
  NOR2X2 \ctrl/add_1_root_add_16_2/U41  ( .A(n513), .B(mux_out[3]), .Y(
        \ctrl/add_1_root_add_16_2/n36 ) );
  NOR2X1 \round/r298/U62  ( .A(\round/r298/n64 ), .B(\round/r298/n52 ), .Y(
        \round/r298/n51 ) );
  OAI21X1 \ctrl/add_1_root_add_16_2/U14  ( .A0(\ctrl/add_1_root_add_16_2/n24 ), 
        .A1(\ctrl/add_1_root_add_16_2/n18 ), .B0(
        \ctrl/add_1_root_add_16_2/n19 ), .Y(\ctrl/add_1_root_add_16_2/n17 ) );
  NOR2X2 \mul/mult_6/U1205  ( .A(sig_B[12]), .B(sig_B[13]), .Y(
        \mul/mult_6/n644 ) );
  XNOR2X2 \mul/mult_6/U1058  ( .A(sig_A[17]), .B(sig_A[18]), .Y(
        \mul/mult_6/n1437 ) );
  NOR2X2 \mul/mult_6/U1299  ( .A(sig_B[1]), .B(sig_B[2]), .Y(\mul/mult_6/n705 ) );
  NOR2X2 \mul/mult_6/U1293  ( .A(sig_B[2]), .B(sig_B[3]), .Y(\mul/mult_6/n702 ) );
  XNOR2X1 \mul/mult_6/U1099  ( .A(sig_A[0]), .B(sig_A[1]), .Y(
        \mul/mult_6/n1451 ) );
  NOR2X2 \mul/mult_6/U1276  ( .A(sig_B[4]), .B(sig_B[5]), .Y(\mul/mult_6/n691 ) );
  XNOR2X2 \mul/mult_6/U1051  ( .A(sig_A[20]), .B(sig_A[21]), .Y(
        \mul/mult_6/n1436 ) );
  NOR2X2 \mul/mult_6/U1251  ( .A(sig_B[7]), .B(sig_B[8]), .Y(\mul/mult_6/n675 ) );
  NOR2X2 \mul/mult_6/U1185  ( .A(sig_B[14]), .B(sig_B[15]), .Y(
        \mul/mult_6/n630 ) );
  NOR2X2 \mul/mult_6/U1146  ( .A(sig_B[18]), .B(sig_B[19]), .Y(
        \mul/mult_6/n603 ) );
  NOR2X2 \mul/mult_6/U1128  ( .A(sig_B[20]), .B(sig_B[21]), .Y(
        \mul/mult_6/n591 ) );
  ADDFX1 \expadd/add_0_root_sub_0_root_sub_8/U6  ( .A(\expadd/N3 ), .B(
        exp_B[3]), .CI(\expadd/add_0_root_sub_0_root_sub_8/n7 ), .CO(
        \expadd/add_0_root_sub_0_root_sub_8/n6 ), .S(exp_P[3]) );
  OAI21XL \mul/mult_6/U483  ( .A0(n545), .A1(\mul/mult_6/n68 ), .B0(
        \mul/mult_6/n1046 ), .Y(\mul/mult_6/n1020 ) );
  XOR2XL \mul/mult_6/U633  ( .A(\mul/mult_6/n1119 ), .B(sig_A[14]), .Y(
        \mul/mult_6/n829 ) );
  XOR2XL \mul/mult_6/U701  ( .A(\mul/mult_6/n1166 ), .B(sig_A[11]), .Y(
        \mul/mult_6/n851 ) );
  MXI2X1 \align/sra_10/U276  ( .A(\align/sra_10/n278 ), .B(\align/sra_10/n279 ), .S0(n507), .Y(\align/sra_10/n224 ) );
  MXI2X1 \align/sra_10/U200  ( .A(\align/sra_10/n250 ), .B(n706), .S0(
        \align/sra_11/SH[1] ), .Y(\align/sra_10/n200 ) );
  AOI21X4 \sigadd/add_9/U273  ( .A0(\sigadd/add_9/n210 ), .A1(n549), .B0(
        \sigadd/add_9/n207 ), .Y(\sigadd/add_9/n205 ) );
  AOI21X4 \sigadd/add_9/U259  ( .A0(\sigadd/add_9/n202 ), .A1(n548), .B0(
        \sigadd/add_9/n199 ), .Y(\sigadd/add_9/n197 ) );
  AOI21X4 \sigadd/add_9/U245  ( .A0(\sigadd/add_9/n194 ), .A1(n547), .B0(
        \sigadd/add_9/n191 ), .Y(\sigadd/add_9/n189 ) );
  AOI21X4 \sigadd/add_9/U203  ( .A0(\sigadd/add_9/n170 ), .A1(n577), .B0(
        \sigadd/add_9/n167 ), .Y(\sigadd/add_9/n165 ) );
  AOI21X4 \sigadd/add_9/U189  ( .A0(\sigadd/add_9/n162 ), .A1(n576), .B0(
        \sigadd/add_9/n159 ), .Y(\sigadd/add_9/n157 ) );
  AOI21X4 \sigadd/add_9/U175  ( .A0(\sigadd/add_9/n154 ), .A1(n575), .B0(
        \sigadd/add_9/n151 ), .Y(\sigadd/add_9/n149 ) );
  AOI21X4 \sigadd/add_9/U161  ( .A0(\sigadd/add_9/n146 ), .A1(n574), .B0(
        \sigadd/add_9/n143 ), .Y(\sigadd/add_9/n141 ) );
  AOI21X4 \sigadd/add_9/U147  ( .A0(\sigadd/add_9/n138 ), .A1(n573), .B0(
        \sigadd/add_9/n135 ), .Y(\sigadd/add_9/n133 ) );
  AOI21X4 \sigadd/add_9/U133  ( .A0(\sigadd/add_9/n130 ), .A1(n599), .B0(
        \sigadd/add_9/n127 ), .Y(\sigadd/add_9/n125 ) );
  AOI21X4 \sigadd/add_9/U119  ( .A0(\sigadd/add_9/n122 ), .A1(n598), .B0(
        \sigadd/add_9/n119 ), .Y(\sigadd/add_9/n117 ) );
  AOI21X4 \sigadd/add_9/U105  ( .A0(\sigadd/add_9/n114 ), .A1(n597), .B0(
        \sigadd/add_9/n111 ), .Y(\sigadd/add_9/n109 ) );
  AOI21X4 \sigadd/add_9/U91  ( .A0(\sigadd/add_9/n106 ), .A1(n596), .B0(
        \sigadd/add_9/n103 ), .Y(\sigadd/add_9/n101 ) );
  AOI21X4 \sigadd/add_9/U77  ( .A0(\sigadd/add_9/n98 ), .A1(n595), .B0(
        \sigadd/add_9/n95 ), .Y(\sigadd/add_9/n93 ) );
  AOI21X4 \sigadd/add_9/U63  ( .A0(\sigadd/add_9/n90 ), .A1(n594), .B0(
        \sigadd/add_9/n87 ), .Y(\sigadd/add_9/n85 ) );
  OAI21X4 \sigadd/add_9/U57  ( .A0(\sigadd/add_9/n85 ), .A1(\sigadd/add_9/n83 ), .B0(\sigadd/add_9/n84 ), .Y(\sigadd/add_9/n82 ) );
  AOI21X4 \sigadd/add_9/U49  ( .A0(\sigadd/add_9/n82 ), .A1(n593), .B0(
        \sigadd/add_9/n79 ), .Y(\sigadd/add_9/n77 ) );
  OAI21X4 \sigadd/add_9/U43  ( .A0(\sigadd/add_9/n77 ), .A1(\sigadd/add_9/n75 ), .B0(\sigadd/add_9/n76 ), .Y(\sigadd/add_9/n74 ) );
  OAI21X4 \sigadd/add_9/U29  ( .A0(\sigadd/add_9/n69 ), .A1(\sigadd/add_9/n67 ), .B0(\sigadd/add_9/n68 ), .Y(\sigadd/add_9/n66 ) );
  NOR2X2 \ctrl/add_1_root_add_16_2/U17  ( .A(n504), .B(mux_out[5]), .Y(
        \ctrl/add_1_root_add_16_2/n18 ) );
  NOR2X1 \normal/sll_15/U46  ( .A(\normal/sll_15/n1 ), .B(n503), .Y(
        \normal/N49 ) );
  NAND2X2 \round/r298/U40  ( .A(norm_out[21]), .B(norm_out[20]), .Y(
        \round/r298/n31 ) );
  NAND2XL \round/r298/U57  ( .A(\round/r298/n53 ), .B(norm_out[18]), .Y(
        \round/r298/n47 ) );
  NAND2XL \round/r298/U75  ( .A(\round/r298/n84 ), .B(\round/r298/n63 ), .Y(
        \round/r298/n62 ) );
  OAI21X1 \mul/mult_6/U1273  ( .A0(\mul/mult_6/n691 ), .A1(\mul/mult_6/n697 ), 
        .B0(\mul/mult_6/n692 ), .Y(\mul/mult_6/n690 ) );
  XNOR2X2 \mul/mult_6/U1079  ( .A(sig_A[8]), .B(sig_A[9]), .Y(
        \mul/mult_6/n1440 ) );
  NAND2X2 \mul/mult_6/U1307  ( .A(sig_B[0]), .B(sig_B[1]), .Y(
        \mul/mult_6/n707 ) );
  NOR2X2 \mul/mult_6/U1262  ( .A(sig_B[6]), .B(sig_B[7]), .Y(\mul/mult_6/n683 ) );
  XNOR2X2 \mul/mult_6/U1086  ( .A(sig_A[5]), .B(sig_A[6]), .Y(
        \mul/mult_6/n1441 ) );
  NOR2X2 \mul/mult_6/U1245  ( .A(sig_B[8]), .B(sig_B[9]), .Y(\mul/mult_6/n672 ) );
  XNOR2X2 \mul/mult_6/U1065  ( .A(sig_A[14]), .B(sig_A[15]), .Y(
        \mul/mult_6/n1438 ) );
  OAI21X1 \mul/mult_6/U1161  ( .A0(\mul/mult_6/n615 ), .A1(\mul/mult_6/n621 ), 
        .B0(\mul/mult_6/n616 ), .Y(\mul/mult_6/n614 ) );
  OAI21X1 \mul/mult_6/U1242  ( .A0(\mul/mult_6/n672 ), .A1(\mul/mult_6/n676 ), 
        .B0(\mul/mult_6/n673 ), .Y(\mul/mult_6/n671 ) );
  AOI21X1 \mul/mult_6/U1141  ( .A0(\mul/mult_6/n601 ), .A1(\mul/mult_6/n614 ), 
        .B0(\mul/mult_6/n602 ), .Y(\mul/mult_6/n600 ) );
  OAI21X1 \mul/mult_6/U990  ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n8 ), 
        .B0(n523), .Y(\mul/mult_6/n1335 ) );
  OAI21X1 \mul/mult_6/U987  ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n8 ), 
        .B0(\mul/mult_6/n1360 ), .Y(\mul/mult_6/n1334 ) );
  AOI21X1 \mul/mult_6/U1271  ( .A0(\mul/mult_6/n698 ), .A1(\mul/mult_6/n689 ), 
        .B0(\mul/mult_6/n690 ), .Y(\mul/mult_6/n688 ) );
  OAI21X1 \mul/mult_6/U1196  ( .A0(\mul/mult_6/n677 ), .A1(\mul/mult_6/n638 ), 
        .B0(\mul/mult_6/n639 ), .Y(\mul/mult_6/n637 ) );
  OAI21X1 \mul/mult_6/U1157  ( .A0(\mul/mult_6/n623 ), .A1(\mul/mult_6/n611 ), 
        .B0(\mul/mult_6/n612 ), .Y(\mul/mult_6/n610 ) );
  ADDFXL \mul/mult_6/U195  ( .A(sig_B[16]), .B(n672), .CI(\mul/mult_6/n786 ), 
        .CO(\mul/mult_6/n205 ), .S(\mul/mult_6/n206 ) );
  CLKNAND2X2 \sigadd/add_9/U2  ( .A(n539), .B(\sigadd/add_9/n52 ), .Y(
        \sigadd/add_9/n1 ) );
  OAI21X4 \sigadd/add_9/U295  ( .A0(\sigadd/add_9/n221 ), .A1(
        \sigadd/add_9/n219 ), .B0(\sigadd/add_9/n220 ), .Y(\sigadd/add_9/n218 ) );
  OAI21X4 \sigadd/add_9/U281  ( .A0(\sigadd/add_9/n213 ), .A1(
        \sigadd/add_9/n211 ), .B0(\sigadd/add_9/n212 ), .Y(\sigadd/add_9/n210 ) );
  OAI21X4 \sigadd/add_9/U267  ( .A0(\sigadd/add_9/n205 ), .A1(
        \sigadd/add_9/n203 ), .B0(\sigadd/add_9/n204 ), .Y(\sigadd/add_9/n202 ) );
  AOI21X4 \sigadd/add_9/U7  ( .A0(\sigadd/add_9/n58 ), .A1(n617), .B0(
        \sigadd/add_9/n55 ), .Y(\sigadd/add_9/n53 ) );
  CLKNAND2X2 \ctrl/add_1_root_add_16_2/U65  ( .A(n534), .B(
        \ctrl/add_1_root_add_16_2/n57 ), .Y(\ctrl/add_1_root_add_16_2/n5 ) );
  AOI21X1 \ctrl/add_1_root_add_16_2/U24  ( .A0(\ctrl/add_1_root_add_16_2/n31 ), 
        .A1(n533), .B0(\ctrl/add_1_root_add_16_2/n26 ), .Y(
        \ctrl/add_1_root_add_16_2/n24 ) );
  NOR2X2 \ctrl/sub_0_root_add_0_root_sub_16/U31  ( .A(
        \ctrl/sub_0_root_add_0_root_sub_16/A[3] ), .B(n709), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n25 ) );
  CLKXOR2X2 U653 ( .A(\sigadd/add_9/n49 ), .B(\sigadd/add_9/n246 ), .Y(
        \sigadd/sig[1] ) );
  NOR2X4 U654 ( .A(\round/r298/n113 ), .B(\round/r298/n106 ), .Y(
        \round/r298/n105 ) );
  OAI22X1 U655 ( .A0(n881), .A1(n880), .B0(n884), .B1(n942), .Y(n937) );
  INVX2 U656 ( .A(\round/r298/n85 ), .Y(\round/r298/n84 ) );
  MX2X1 U657 ( .A(\normal/N26 ), .B(\normal/N72 ), .S0(n999), .Y(norm_out[4])
         );
  MX2X1 U658 ( .A(\normal/N28 ), .B(\normal/N74 ), .S0(n999), .Y(norm_out[6])
         );
  MX2X1 U659 ( .A(\normal/N30 ), .B(\normal/N76 ), .S0(n999), .Y(norm_out[8])
         );
  MX2X1 U660 ( .A(\normal/N31 ), .B(\normal/N77 ), .S0(n999), .Y(norm_out[9])
         );
  MX2X1 U661 ( .A(\normal/N42 ), .B(\normal/N88 ), .S0(n999), .Y(norm_out[20])
         );
  MXI2X1 U662 ( .A(\normal/srl_15/n72 ), .B(\normal/srl_15/n76 ), .S0(n512), 
        .Y(\normal/srl_15/n24 ) );
  NAND3XL U663 ( .A(n986), .B(n985), .C(n984), .Y(zero_cnt[0]) );
  NAND3XL U664 ( .A(n935), .B(n934), .C(n933), .Y(n936) );
  NAND2X4 U665 ( .A(n1039), .B(mux_out[3]), .Y(n1038) );
  NOR2X2 U666 ( .A(\round/r298/n31 ), .B(\round/r298/n21 ), .Y(
        \round/r298/n18 ) );
  NAND2X2 U667 ( .A(\round/r298/n86 ), .B(\round/r298/n105 ), .Y(
        \round/r298/n85 ) );
  NAND2X2 U668 ( .A(n1036), .B(mux_out[5]), .Y(n1035) );
  MX2X1 U669 ( .A(\normal/N43 ), .B(\normal/N89 ), .S0(n999), .Y(norm_out[21])
         );
  NOR2X2 U670 ( .A(n704), .B(\ctrl/add_1_root_add_16_2/A[2] ), .Y(
        \ctrl/add_1_root_add_16_2/n41 ) );
  NAND2X2 U671 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/A[5] ), .B(n713), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n14 ) );
  BUFX2 U672 ( .A(n39), .Y(n702) );
  INVX4 U673 ( .A(\sigadd/sub_add_11_b0/B[49] ), .Y(n661) );
  OAI211XL U674 ( .A0(n522), .A1(n1007), .B0(n1006), .C0(n1005), .Y(D[0]) );
  AOI222XL U675 ( .A0(norm_out[4]), .A1(n1026), .B0(\round/N9 ), .B1(n662), 
        .C0(n39), .C1(\round/N10 ), .Y(n1008) );
  AOI222XL U676 ( .A0(norm_out[5]), .A1(n1026), .B0(n662), .B1(\round/N10 ), 
        .C0(n39), .C1(\round/N11 ), .Y(n1009) );
  AOI222XL U677 ( .A0(norm_out[6]), .A1(n1026), .B0(n662), .B1(\round/N11 ), 
        .C0(n39), .C1(\round/N12 ), .Y(n1010) );
  AOI222XL U678 ( .A0(norm_out[7]), .A1(n1026), .B0(n1025), .B1(\round/N12 ), 
        .C0(n39), .C1(\round/N13 ), .Y(n1011) );
  AOI222XL U679 ( .A0(norm_out[8]), .A1(n1026), .B0(n1025), .B1(\round/N13 ), 
        .C0(n39), .C1(\round/N14 ), .Y(n1012) );
  AOI222XL U680 ( .A0(norm_out[9]), .A1(n1026), .B0(n662), .B1(\round/N14 ), 
        .C0(n39), .C1(\round/N15 ), .Y(n1013) );
  AOI222XL U681 ( .A0(norm_out[10]), .A1(n1026), .B0(n662), .B1(\round/N15 ), 
        .C0(n39), .C1(\round/N16 ), .Y(n1014) );
  AOI222XL U682 ( .A0(norm_out[11]), .A1(n1026), .B0(n1025), .B1(\round/N16 ), 
        .C0(n39), .C1(\round/N17 ), .Y(n1015) );
  AOI222XL U683 ( .A0(norm_out[12]), .A1(n1026), .B0(n1025), .B1(\round/N17 ), 
        .C0(n39), .C1(\round/N18 ), .Y(n1016) );
  AOI222XL U684 ( .A0(norm_out[13]), .A1(n1026), .B0(n662), .B1(\round/N18 ), 
        .C0(n39), .C1(\round/N19 ), .Y(n1017) );
  AOI222XL U685 ( .A0(norm_out[14]), .A1(n1026), .B0(n662), .B1(\round/N19 ), 
        .C0(n39), .C1(\round/N20 ), .Y(n1018) );
  AOI222XL U686 ( .A0(norm_out[15]), .A1(n1026), .B0(n1025), .B1(\round/N20 ), 
        .C0(n39), .C1(\round/N21 ), .Y(n1019) );
  AOI222XL U687 ( .A0(norm_out[16]), .A1(n1026), .B0(n1025), .B1(\round/N21 ), 
        .C0(n39), .C1(\round/N22 ), .Y(n1020) );
  AOI222XL U688 ( .A0(norm_out[17]), .A1(n1026), .B0(n662), .B1(\round/N22 ), 
        .C0(n39), .C1(\round/N23 ), .Y(n1021) );
  AOI222XL U689 ( .A0(norm_out[18]), .A1(n1026), .B0(n662), .B1(\round/N23 ), 
        .C0(n39), .C1(\round/N24 ), .Y(n1022) );
  AOI222XL U690 ( .A0(norm_out[19]), .A1(n1026), .B0(n1025), .B1(\round/N24 ), 
        .C0(n39), .C1(\round/N25 ), .Y(n1023) );
  AOI222XL U691 ( .A0(norm_out[20]), .A1(n1026), .B0(n1025), .B1(\round/N25 ), 
        .C0(n39), .C1(\round/N26 ), .Y(n1024) );
  INVX8 U692 ( .A(n1043), .Y(n999) );
  CLKBUFX16 U693 ( .A(n1030), .Y(n516) );
  OAI21X2 U694 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n560), .B0(n831), .Y(
        add_out[48]) );
  CLKBUFX4 U695 ( .A(\mul/mult_6/n12 ), .Y(n681) );
  BUFX10 U696 ( .A(n519), .Y(n508) );
  NOR3X1 U697 ( .A(\normal/srl_15/A[36] ), .B(add_out[35]), .C(add_out[34]), 
        .Y(n836) );
  OAI21X1 U698 ( .A0(\mul/mult_6/n699 ), .A1(\mul/mult_6/n679 ), .B0(
        \mul/mult_6/n680 ), .Y(\mul/mult_6/n678 ) );
  OAI211XL U699 ( .A0(add_out[19]), .A1(add_out[20]), .B0(n875), .C0(n871), 
        .Y(n955) );
  XNOR2X2 U700 ( .A(sig_A[2]), .B(sig_A[3]), .Y(\mul/mult_6/n1442 ) );
  MXI2X1 U701 ( .A(\align/sra_10/n222 ), .B(\align/sra_10/n224 ), .S0(
        \align/sra_11/SH[1] ), .Y(\align/sra_10/n172 ) );
  OAI211XL U702 ( .A0(n940), .A1(n873), .B0(n872), .C0(n955), .Y(n892) );
  OAI211XL U703 ( .A0(n970), .A1(n956), .B0(n885), .C0(n870), .Y(n959) );
  OAI21X1 U704 ( .A0(\mul/mult_6/n677 ), .A1(\mul/mult_6/n652 ), .B0(
        \mul/mult_6/n653 ), .Y(\mul/mult_6/n651 ) );
  MXI2X1 U705 ( .A(\align/sra_10/n192 ), .B(\align/sra_10/n196 ), .S0(n505), 
        .Y(\align/sra_10/n142 ) );
  OAI21X1 U706 ( .A0(\mul/mult_6/n677 ), .A1(\mul/mult_6/n668 ), .B0(
        \mul/mult_6/n669 ), .Y(\mul/mult_6/n667 ) );
  MXI2X1 U707 ( .A(\align/sra_10/n176 ), .B(\align/sra_10/n180 ), .S0(n511), 
        .Y(\align/sra_10/n126 ) );
  MXI2X1 U708 ( .A(\align/sra_10/n184 ), .B(\align/sra_10/n188 ), .S0(n511), 
        .Y(\align/sra_10/n134 ) );
  OAI21X1 U709 ( .A0(n502), .A1(n557), .B0(n727), .Y(sel_P[48]) );
  OAI21X1 U710 ( .A0(n886), .A1(n942), .B0(n885), .Y(n915) );
  OAI31X1 U711 ( .A0(n964), .A1(n963), .A2(\normal/srl_15/A[9] ), .B0(n962), 
        .Y(n965) );
  AOI21X1 U712 ( .A0(\mul/mult_6/n700 ), .A1(\mul/mult_6/n708 ), .B0(
        \mul/mult_6/n701 ), .Y(\mul/mult_6/n699 ) );
  NOR2X2 U713 ( .A(\mul/mult_6/n1439 ), .B(\mul/mult_6/n1455 ), .Y(
        \mul/mult_6/n42 ) );
  AOI21X1 U714 ( .A0(n901), .A1(n900), .B0(n899), .Y(n985) );
  AOI222XL U715 ( .A0(n681), .A1(sig_B[6]), .B0(\mul/mult_6/n543 ), .B1(
        sig_B[5]), .C0(\mul/mult_6/n20 ), .C1(sig_B[4]), .Y(\mul/mult_6/n1304 ) );
  AOI222XL U716 ( .A0(n681), .A1(sig_B[4]), .B0(n700), .B1(sig_B[3]), .C0(
        \mul/mult_6/n20 ), .C1(sig_B[2]), .Y(\mul/mult_6/n1306 ) );
  AOI222XL U717 ( .A0(n683), .A1(sig_B[4]), .B0(n699), .B1(sig_B[3]), .C0(
        \mul/mult_6/n30 ), .C1(sig_B[2]), .Y(\mul/mult_6/n1254 ) );
  AOI222XL U718 ( .A0(n679), .A1(sig_B[2]), .B0(n701), .B1(sig_B[1]), .C0(
        \mul/mult_6/n9 ), .C1(sig_B[0]), .Y(\mul/mult_6/n1360 ) );
  AOI222XL U719 ( .A0(n681), .A1(sig_B[3]), .B0(n700), .B1(sig_B[2]), .C0(
        \mul/mult_6/n20 ), .C1(sig_B[1]), .Y(\mul/mult_6/n1307 ) );
  AOI222XL U720 ( .A0(n681), .A1(sig_B[2]), .B0(n700), .B1(sig_B[1]), .C0(
        \mul/mult_6/n20 ), .C1(sig_B[0]), .Y(\mul/mult_6/n1308 ) );
  AOI222XL U721 ( .A0(n683), .A1(sig_B[3]), .B0(n699), .B1(sig_B[2]), .C0(
        \mul/mult_6/n30 ), .C1(sig_B[1]), .Y(\mul/mult_6/n1255 ) );
  AOI222XL U722 ( .A0(n683), .A1(sig_B[2]), .B0(n699), .B1(sig_B[1]), .C0(
        \mul/mult_6/n30 ), .C1(sig_B[0]), .Y(\mul/mult_6/n1256 ) );
  AOI222XL U723 ( .A0(n685), .A1(sig_B[3]), .B0(n698), .B1(sig_B[2]), .C0(
        \mul/mult_6/n40 ), .C1(sig_B[1]), .Y(\mul/mult_6/n1203 ) );
  AOI222XL U724 ( .A0(n685), .A1(sig_B[2]), .B0(n698), .B1(sig_B[1]), .C0(
        \mul/mult_6/n40 ), .C1(sig_B[0]), .Y(\mul/mult_6/n1204 ) );
  AOI222XL U725 ( .A0(n679), .A1(sig_B[4]), .B0(n701), .B1(sig_B[3]), .C0(
        \mul/mult_6/n9 ), .C1(sig_B[2]), .Y(\mul/mult_6/n1358 ) );
  AOI222XL U726 ( .A0(n679), .A1(sig_B[5]), .B0(n701), .B1(sig_B[4]), .C0(
        \mul/mult_6/n9 ), .C1(sig_B[3]), .Y(\mul/mult_6/n1357 ) );
  AOI222XL U727 ( .A0(n679), .A1(sig_B[6]), .B0(n701), .B1(sig_B[5]), .C0(
        \mul/mult_6/n9 ), .C1(sig_B[4]), .Y(\mul/mult_6/n1356 ) );
  AOI222XL U728 ( .A0(n679), .A1(sig_B[8]), .B0(\mul/mult_6/n547 ), .B1(
        sig_B[7]), .C0(\mul/mult_6/n9 ), .C1(sig_B[6]), .Y(\mul/mult_6/n1354 )
         );
  AOI222XL U729 ( .A0(n679), .A1(sig_B[3]), .B0(n701), .B1(sig_B[2]), .C0(
        \mul/mult_6/n9 ), .C1(sig_B[1]), .Y(\mul/mult_6/n1359 ) );
  NOR2X2 U730 ( .A(\mul/mult_6/n1441 ), .B(\mul/mult_6/n1457 ), .Y(
        \mul/mult_6/n22 ) );
  NOR2X2 U731 ( .A(\mul/mult_6/n1440 ), .B(\mul/mult_6/n1456 ), .Y(
        \mul/mult_6/n32 ) );
  NAND2X2 U732 ( .A(n562), .B(\mul/mult_6/n707 ), .Y(\mul/mult_6/n1387 ) );
  CLKXOR2X2 U733 ( .A(\mul/mult_6/n651 ), .B(\mul/mult_6/n562 ), .Y(n572) );
  CLKXOR2X2 U734 ( .A(\mul/mult_6/n667 ), .B(\mul/mult_6/n564 ), .Y(n542) );
  CLKXOR2X2 U735 ( .A(\mul/mult_6/n674 ), .B(\mul/mult_6/n565 ), .Y(n543) );
  CLKXOR2X2 U736 ( .A(\mul/mult_6/n704 ), .B(\mul/mult_6/n571 ), .Y(n546) );
  CLKXOR2X2 U737 ( .A(\mul/mult_6/n685 ), .B(\mul/mult_6/n567 ), .Y(n544) );
  INVX2 U738 ( .A(\mul/mult_6/n1407 ), .Y(\mul/mult_6/n1382 ) );
  INVX2 U739 ( .A(\mul/mult_6/n1411 ), .Y(\mul/mult_6/n1386 ) );
  INVX2 U740 ( .A(\mul/mult_6/n1402 ), .Y(\mul/mult_6/n1377 ) );
  INVX2 U741 ( .A(\mul/mult_6/n1400 ), .Y(\mul/mult_6/n1375 ) );
  INVX2 U742 ( .A(\mul/mult_6/n1408 ), .Y(\mul/mult_6/n1383 ) );
  INVX2 U743 ( .A(\mul/mult_6/n1405 ), .Y(\mul/mult_6/n1380 ) );
  OAI211XL U744 ( .A0(n957), .A1(n956), .B0(n955), .C0(n954), .Y(n958) );
  OAI211XL U745 ( .A0(n878), .A1(n877), .B0(n896), .C0(n876), .Y(n879) );
  OAI211XL U746 ( .A0(n904), .A1(n903), .B0(n902), .C0(n985), .Y(n905) );
  AOI22XL U747 ( .A0(n698), .A1(sig_B[0]), .B0(n685), .B1(sig_B[1]), .Y(n528)
         );
  INVX2 U748 ( .A(\mul/mult_6/n678 ), .Y(\mul/mult_6/n677 ) );
  INVX2 U749 ( .A(sig_A[0]), .Y(\mul/mult_6/n1443 ) );
  XOR2X2 U750 ( .A(sig_A[1]), .B(sig_A[2]), .Y(\mul/mult_6/n1459 ) );
  OR2X2 U751 ( .A(\mul/mult_6/n127 ), .B(sig_B[21]), .Y(\mul/mult_6/n126 ) );
  INVX2 U752 ( .A(sig_P[47]), .Y(\selc/r299/A[47] ) );
  BUFX5 U753 ( .A(\mul/mult_6/n531 ), .Y(n518) );
  CLKBUFX4 U754 ( .A(\mul/mult_6/n62 ), .Y(n692) );
  OAI21X1 U755 ( .A0(\mul/mult_6/n623 ), .A1(\mul/mult_6/n599 ), .B0(
        \mul/mult_6/n600 ), .Y(\mul/mult_6/n598 ) );
  AOI21X1 U756 ( .A0(\mul/mult_6/n658 ), .A1(\mul/mult_6/n671 ), .B0(
        \mul/mult_6/n659 ), .Y(\mul/mult_6/n653 ) );
  AOI21X2 U757 ( .A0(\mul/mult_6/n678 ), .A1(\mul/mult_6/n624 ), .B0(
        \mul/mult_6/n625 ), .Y(\mul/mult_6/n623 ) );
  NOR2X2 U758 ( .A(\mul/mult_6/n1438 ), .B(\mul/mult_6/n1454 ), .Y(
        \mul/mult_6/n52 ) );
  AOI222XL U759 ( .A0(n681), .A1(sig_B[7]), .B0(\mul/mult_6/n543 ), .B1(
        sig_B[6]), .C0(\mul/mult_6/n20 ), .C1(sig_B[5]), .Y(\mul/mult_6/n1303 ) );
  AOI222XL U760 ( .A0(n689), .A1(sig_B[2]), .B0(n690), .B1(sig_B[1]), .C0(
        \mul/mult_6/n60 ), .C1(sig_B[0]), .Y(\mul/mult_6/n1100 ) );
  AOI222XL U761 ( .A0(n692), .A1(sig_B[2]), .B0(n693), .B1(sig_B[1]), .C0(
        \mul/mult_6/n70 ), .C1(sig_B[0]), .Y(\mul/mult_6/n1048 ) );
  AOI222XL U762 ( .A0(n689), .A1(sig_B[4]), .B0(\mul/mult_6/n54 ), .B1(
        sig_B[3]), .C0(\mul/mult_6/n60 ), .C1(sig_B[2]), .Y(\mul/mult_6/n1098 ) );
  AOI222XL U763 ( .A0(n689), .A1(sig_B[3]), .B0(n690), .B1(sig_B[2]), .C0(
        \mul/mult_6/n60 ), .C1(sig_B[1]), .Y(\mul/mult_6/n1099 ) );
  AOI222XL U764 ( .A0(n681), .A1(sig_B[8]), .B0(\mul/mult_6/n543 ), .B1(
        sig_B[7]), .C0(\mul/mult_6/n20 ), .C1(sig_B[6]), .Y(\mul/mult_6/n1302 ) );
  AOI222XL U765 ( .A0(n687), .A1(sig_B[2]), .B0(n518), .B1(sig_B[1]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[0]), .Y(\mul/mult_6/n1152 ) );
  AOI222XL U766 ( .A0(n679), .A1(sig_B[10]), .B0(\mul/mult_6/n547 ), .B1(
        sig_B[9]), .C0(\mul/mult_6/n9 ), .C1(sig_B[8]), .Y(\mul/mult_6/n1352 )
         );
  AOI222XL U767 ( .A0(n685), .A1(sig_B[4]), .B0(n698), .B1(sig_B[3]), .C0(
        \mul/mult_6/n40 ), .C1(sig_B[2]), .Y(\mul/mult_6/n1202 ) );
  AOI222XL U768 ( .A0(n679), .A1(sig_B[9]), .B0(\mul/mult_6/n547 ), .B1(
        sig_B[8]), .C0(\mul/mult_6/n9 ), .C1(sig_B[7]), .Y(\mul/mult_6/n1353 )
         );
  AOI222XL U769 ( .A0(n687), .A1(sig_B[3]), .B0(n518), .B1(sig_B[2]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[1]), .Y(\mul/mult_6/n1151 ) );
  AOI222XL U770 ( .A0(n687), .A1(sig_B[6]), .B0(n518), .B1(sig_B[5]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[4]), .Y(\mul/mult_6/n1148 ) );
  AOI222XL U771 ( .A0(n687), .A1(sig_B[5]), .B0(n518), .B1(sig_B[4]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[3]), .Y(\mul/mult_6/n1149 ) );
  AOI222XL U772 ( .A0(n687), .A1(sig_B[4]), .B0(n518), .B1(sig_B[3]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[2]), .Y(\mul/mult_6/n1150 ) );
  CLKXOR2X2 U773 ( .A(\mul/mult_6/n598 ), .B(\mul/mult_6/n554 ), .Y(n591) );
  CLKXOR2X2 U774 ( .A(\mul/mult_6/n610 ), .B(\mul/mult_6/n556 ), .Y(n569) );
  CLKXOR2X2 U775 ( .A(\mul/mult_6/n637 ), .B(\mul/mult_6/n560 ), .Y(n571) );
  CLKXOR2X2 U776 ( .A(\mul/mult_6/n622 ), .B(\mul/mult_6/n558 ), .Y(n570) );
  INVX2 U777 ( .A(\mul/mult_6/n1391 ), .Y(\mul/mult_6/n1366 ) );
  INVX2 U778 ( .A(\mul/mult_6/n1390 ), .Y(\mul/mult_6/n1365 ) );
  INVX2 U779 ( .A(\mul/mult_6/n1396 ), .Y(\mul/mult_6/n1371 ) );
  INVX2 U780 ( .A(\mul/mult_6/n1392 ), .Y(\mul/mult_6/n1367 ) );
  INVX2 U781 ( .A(\mul/mult_6/n1394 ), .Y(\mul/mult_6/n1369 ) );
  INVX2 U782 ( .A(\mul/mult_6/n1398 ), .Y(\mul/mult_6/n1373 ) );
  AOI22XL U783 ( .A0(n693), .A1(sig_B[0]), .B0(n692), .B1(sig_B[1]), .Y(n610)
         );
  AOI22XL U784 ( .A0(n518), .A1(sig_B[0]), .B0(n687), .B1(sig_B[1]), .Y(n527)
         );
  AOI22XL U785 ( .A0(n690), .A1(sig_B[0]), .B0(n689), .B1(sig_B[1]), .Y(n535)
         );
  CLKBUFX4 U786 ( .A(\mul/mult_6/n74 ), .Y(n696) );
  AOI222XL U787 ( .A0(n683), .A1(sig_B[14]), .B0(\mul/mult_6/n539 ), .B1(
        sig_B[13]), .C0(\mul/mult_6/n30 ), .C1(sig_B[12]), .Y(
        \mul/mult_6/n1244 ) );
  AOI222XL U788 ( .A0(n689), .A1(sig_B[5]), .B0(\mul/mult_6/n54 ), .B1(
        sig_B[4]), .C0(\mul/mult_6/n60 ), .C1(sig_B[3]), .Y(\mul/mult_6/n1097 ) );
  AOI222XL U789 ( .A0(n689), .A1(sig_B[11]), .B0(n690), .B1(sig_B[10]), .C0(
        \mul/mult_6/n60 ), .C1(sig_B[9]), .Y(\mul/mult_6/n1091 ) );
  AOI222XL U790 ( .A0(n692), .A1(sig_B[8]), .B0(n693), .B1(sig_B[7]), .C0(
        \mul/mult_6/n70 ), .C1(sig_B[6]), .Y(\mul/mult_6/n1042 ) );
  AOI222XL U791 ( .A0(n685), .A1(sig_B[18]), .B0(n698), .B1(sig_B[17]), .C0(
        \mul/mult_6/n40 ), .C1(sig_B[16]), .Y(\mul/mult_6/n1188 ) );
  AOI222XL U792 ( .A0(n692), .A1(sig_B[10]), .B0(n693), .B1(sig_B[9]), .C0(
        \mul/mult_6/n70 ), .C1(sig_B[8]), .Y(\mul/mult_6/n1040 ) );
  AOI222XL U793 ( .A0(n692), .A1(sig_B[3]), .B0(n693), .B1(sig_B[2]), .C0(
        \mul/mult_6/n70 ), .C1(sig_B[1]), .Y(\mul/mult_6/n1047 ) );
  AOI222XL U794 ( .A0(n689), .A1(sig_B[12]), .B0(n690), .B1(sig_B[11]), .C0(
        \mul/mult_6/n60 ), .C1(sig_B[10]), .Y(\mul/mult_6/n1090 ) );
  AOI222XL U795 ( .A0(n692), .A1(sig_B[4]), .B0(n693), .B1(sig_B[3]), .C0(
        \mul/mult_6/n70 ), .C1(sig_B[2]), .Y(\mul/mult_6/n1046 ) );
  AOI222XL U796 ( .A0(n695), .A1(sig_B[3]), .B0(n696), .B1(sig_B[2]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[1]), .Y(\mul/mult_6/n995 ) );
  AOI222XL U797 ( .A0(n695), .A1(sig_B[7]), .B0(n696), .B1(sig_B[6]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[5]), .Y(\mul/mult_6/n991 ) );
  AOI222XL U798 ( .A0(n695), .A1(sig_B[4]), .B0(n696), .B1(sig_B[3]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[2]), .Y(\mul/mult_6/n994 ) );
  INVX2 U799 ( .A(\mul/mult_6/n1364 ), .Y(\mul/mult_6/n1363 ) );
  AOI22XL U800 ( .A0(n696), .A1(sig_B[0]), .B0(n695), .B1(sig_B[1]), .Y(n538)
         );
  AOI222XL U801 ( .A0(n692), .A1(sig_B[16]), .B0(\mul/mult_6/n64 ), .B1(
        sig_B[15]), .C0(\mul/mult_6/n70 ), .C1(sig_B[14]), .Y(
        \mul/mult_6/n1034 ) );
  AOI222XL U802 ( .A0(\mul/mult_6/n42 ), .A1(sig_B[21]), .B0(n518), .B1(
        sig_B[20]), .C0(\mul/mult_6/n50 ), .C1(sig_B[19]), .Y(
        \mul/mult_6/n1133 ) );
  AOI222XL U803 ( .A0(\mul/mult_6/n42 ), .A1(sig_B[20]), .B0(n518), .B1(
        sig_B[19]), .C0(\mul/mult_6/n50 ), .C1(sig_B[18]), .Y(
        \mul/mult_6/n1134 ) );
  AOI222XL U804 ( .A0(n687), .A1(sig_B[17]), .B0(n518), .B1(sig_B[16]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[15]), .Y(\mul/mult_6/n1137 ) );
  AOI222XL U805 ( .A0(n687), .A1(sig_B[18]), .B0(n518), .B1(sig_B[17]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[16]), .Y(\mul/mult_6/n1136 ) );
  AOI222XL U806 ( .A0(n687), .A1(sig_B[16]), .B0(n518), .B1(sig_B[15]), .C0(
        \mul/mult_6/n50 ), .C1(sig_B[14]), .Y(\mul/mult_6/n1138 ) );
  AOI222XL U807 ( .A0(n689), .A1(sig_B[18]), .B0(\mul/mult_6/n54 ), .B1(
        sig_B[17]), .C0(\mul/mult_6/n60 ), .C1(sig_B[16]), .Y(
        \mul/mult_6/n1084 ) );
  AOI222XL U808 ( .A0(n692), .A1(sig_B[11]), .B0(n693), .B1(sig_B[10]), .C0(
        \mul/mult_6/n70 ), .C1(sig_B[9]), .Y(\mul/mult_6/n1039 ) );
  AOI222XL U809 ( .A0(n689), .A1(sig_B[15]), .B0(\mul/mult_6/n54 ), .B1(
        sig_B[14]), .C0(\mul/mult_6/n60 ), .C1(sig_B[13]), .Y(
        \mul/mult_6/n1087 ) );
  AOI222XL U810 ( .A0(n692), .A1(sig_B[13]), .B0(n693), .B1(sig_B[12]), .C0(
        \mul/mult_6/n70 ), .C1(sig_B[11]), .Y(\mul/mult_6/n1037 ) );
  AOI222XL U811 ( .A0(n695), .A1(sig_B[8]), .B0(n696), .B1(sig_B[7]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[6]), .Y(\mul/mult_6/n990 ) );
  AOI222XL U812 ( .A0(n695), .A1(sig_B[9]), .B0(n696), .B1(sig_B[8]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[7]), .Y(\mul/mult_6/n989 ) );
  AOI222XL U813 ( .A0(n695), .A1(sig_B[10]), .B0(n696), .B1(sig_B[9]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[8]), .Y(\mul/mult_6/n988 ) );
  AOI222XL U814 ( .A0(n695), .A1(sig_B[13]), .B0(n696), .B1(sig_B[12]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[11]), .Y(\mul/mult_6/n985 ) );
  AOI222XL U815 ( .A0(n695), .A1(sig_B[12]), .B0(n696), .B1(sig_B[11]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[10]), .Y(\mul/mult_6/n986 ) );
  AOI222XL U816 ( .A0(n695), .A1(sig_B[14]), .B0(n696), .B1(sig_B[13]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[12]), .Y(\mul/mult_6/n984 ) );
  CLKBUFX16 U817 ( .A(sub_out[5]), .Y(n515) );
  AOI222XL U818 ( .A0(\mul/mult_6/n42 ), .A1(sig_B[22]), .B0(n518), .B1(
        sig_B[21]), .C0(\mul/mult_6/n50 ), .C1(sig_B[20]), .Y(
        \mul/mult_6/n1132 ) );
  AOI222XL U819 ( .A0(n692), .A1(sig_B[17]), .B0(\mul/mult_6/n64 ), .B1(
        sig_B[16]), .C0(\mul/mult_6/n70 ), .C1(sig_B[15]), .Y(
        \mul/mult_6/n1033 ) );
  AOI222XL U820 ( .A0(n689), .A1(sig_B[19]), .B0(\mul/mult_6/n54 ), .B1(
        sig_B[18]), .C0(\mul/mult_6/n60 ), .C1(sig_B[17]), .Y(
        \mul/mult_6/n1083 ) );
  AOI222XL U821 ( .A0(\mul/mult_6/n62 ), .A1(sig_B[18]), .B0(\mul/mult_6/n64 ), 
        .B1(sig_B[17]), .C0(\mul/mult_6/n70 ), .C1(sig_B[16]), .Y(
        \mul/mult_6/n1032 ) );
  AOI222XL U822 ( .A0(\mul/mult_6/n62 ), .A1(sig_B[20]), .B0(\mul/mult_6/n64 ), 
        .B1(sig_B[19]), .C0(\mul/mult_6/n70 ), .C1(sig_B[18]), .Y(
        \mul/mult_6/n1030 ) );
  AOI222XL U823 ( .A0(\mul/mult_6/n52 ), .A1(sig_B[22]), .B0(\mul/mult_6/n54 ), 
        .B1(sig_B[21]), .C0(\mul/mult_6/n60 ), .C1(sig_B[20]), .Y(
        \mul/mult_6/n1080 ) );
  AOI222XL U824 ( .A0(\mul/mult_6/n62 ), .A1(sig_B[19]), .B0(\mul/mult_6/n64 ), 
        .B1(sig_B[18]), .C0(\mul/mult_6/n70 ), .C1(sig_B[17]), .Y(
        \mul/mult_6/n1031 ) );
  AOI222XL U825 ( .A0(\mul/mult_6/n62 ), .A1(sig_B[22]), .B0(\mul/mult_6/n64 ), 
        .B1(sig_B[21]), .C0(\mul/mult_6/n70 ), .C1(sig_B[20]), .Y(
        \mul/mult_6/n1028 ) );
  AOI222XL U826 ( .A0(\mul/mult_6/n52 ), .A1(sig_B[21]), .B0(\mul/mult_6/n54 ), 
        .B1(sig_B[20]), .C0(\mul/mult_6/n60 ), .C1(sig_B[19]), .Y(
        \mul/mult_6/n1081 ) );
  AOI222XL U827 ( .A0(\mul/mult_6/n62 ), .A1(sig_B[21]), .B0(\mul/mult_6/n64 ), 
        .B1(sig_B[20]), .C0(\mul/mult_6/n70 ), .C1(sig_B[19]), .Y(
        \mul/mult_6/n1029 ) );
  AOI222XL U828 ( .A0(n695), .A1(sig_B[15]), .B0(n696), .B1(sig_B[14]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[13]), .Y(\mul/mult_6/n983 ) );
  AOI222XL U829 ( .A0(n695), .A1(sig_B[18]), .B0(\mul/mult_6/n74 ), .B1(
        sig_B[17]), .C0(\mul/mult_6/n78 ), .C1(sig_B[16]), .Y(
        \mul/mult_6/n980 ) );
  AOI222XL U830 ( .A0(n695), .A1(sig_B[16]), .B0(n696), .B1(sig_B[15]), .C0(
        \mul/mult_6/n78 ), .C1(sig_B[14]), .Y(\mul/mult_6/n982 ) );
  AOI222XL U831 ( .A0(n695), .A1(sig_B[19]), .B0(\mul/mult_6/n74 ), .B1(
        sig_B[18]), .C0(\mul/mult_6/n78 ), .C1(sig_B[17]), .Y(
        \mul/mult_6/n979 ) );
  AOI222XL U832 ( .A0(n695), .A1(sig_B[20]), .B0(\mul/mult_6/n74 ), .B1(
        sig_B[19]), .C0(\mul/mult_6/n78 ), .C1(sig_B[18]), .Y(
        \mul/mult_6/n978 ) );
  CLKBUFX16 U833 ( .A(n719), .Y(n718) );
  CLKBUFX4 U834 ( .A(n775), .Y(n724) );
  AOI21X1 U835 ( .A0(n514), .A1(\normal/srl_15/n224 ), .B0(n504), .Y(n387) );
  OAI2B1X1 U836 ( .A1N(\normal/srl_15/n222 ), .A0(n514), .B0(n387), .Y(
        \normal/srl_15/n122 ) );
  AOI21X1 U837 ( .A0(n514), .A1(\normal/sll_15/n211 ), .B0(n504), .Y(n388) );
  OAI2B1X1 U838 ( .A1N(\normal/sll_15/n213 ), .A0(n514), .B0(n388), .Y(
        \normal/sll_15/n119 ) );
  AOI21X1 U839 ( .A0(n514), .A1(\normal/sll_15/n216 ), .B0(n504), .Y(n389) );
  OAI2B1X1 U840 ( .A1N(\normal/sll_15/n218 ), .A0(n514), .B0(n389), .Y(
        \normal/sll_15/n124 ) );
  AOI21X1 U841 ( .A0(n514), .A1(\normal/sll_15/n217 ), .B0(n504), .Y(n390) );
  OAI2B1X1 U842 ( .A1N(\normal/sll_15/n219 ), .A0(n514), .B0(n390), .Y(
        \normal/sll_15/n125 ) );
  CLKINVX1 U843 ( .A(n704), .Y(n391) );
  AOI22XL U844 ( .A0(n704), .A1(\normal/sll_15/n50 ), .B0(\normal/sll_15/n54 ), 
        .B1(n391), .Y(n392) );
  AOI22XL U845 ( .A0(n704), .A1(\normal/sll_15/n49 ), .B0(\normal/sll_15/n53 ), 
        .B1(n391), .Y(n393) );
  OAI2B1X1 U846 ( .A1N(n503), .A0(\normal/sll_15/n5 ), .B0(n393), .Y(n394) );
  AOI22XL U847 ( .A0(n704), .A1(\normal/sll_15/n51 ), .B0(\normal/sll_15/n55 ), 
        .B1(n391), .Y(n395) );
  OAI21X1 U848 ( .A0(n503), .A1(\normal/sll_15/n9 ), .B0(n395), .Y(n396) );
  NOR3BX1 U849 ( .AN(n392), .B(n394), .C(n396), .Y(n998) );
  CLKINVX1 U850 ( .A(n503), .Y(n397) );
  AOI22XL U851 ( .A0(n503), .A1(\normal/srl_15/n29 ), .B0(\normal/srl_15/n28 ), 
        .B1(n397), .Y(n398) );
  AOI22XL U852 ( .A0(n503), .A1(\normal/sll_15/n27 ), .B0(\normal/sll_15/n28 ), 
        .B1(n397), .Y(n399) );
  MX2X1 U853 ( .A(n398), .B(n399), .S0(n999), .Y(norm_out[7]) );
  XOR2X1 U854 ( .A(norm_out[20]), .B(\round/r298/n1 ), .Y(\round/N25 ) );
  CLKINVX1 U855 ( .A(n503), .Y(n400) );
  AOI22XL U856 ( .A0(n503), .A1(\normal/srl_15/n46 ), .B0(\normal/srl_15/n45 ), 
        .B1(n400), .Y(n401) );
  AOI22XL U857 ( .A0(n503), .A1(\normal/sll_15/n44 ), .B0(\normal/sll_15/n45 ), 
        .B1(n400), .Y(n402) );
  MX2X1 U858 ( .A(n401), .B(n402), .S0(n999), .Y(norm_out[24]) );
  CLKINVX1 U859 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n10 ), .Y(n403) );
  OAI211X2 U860 ( .A0(\ctrl/sub_0_root_add_0_root_sub_16/n8 ), .A1(
        \ctrl/sub_0_root_add_0_root_sub_16/n19 ), .B0(
        \ctrl/sub_0_root_add_0_root_sub_16/n14 ), .C0(n403), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n7 ) );
  AOI222XL U861 ( .A0(n1026), .A1(norm_out[21]), .B0(n39), .B1(\round/N27 ), 
        .C0(n662), .C1(\round/N26 ), .Y(n404) );
  CLKINVX1 U862 ( .A(n404), .Y(D[18]) );
  OAI2B1X1 U863 ( .A1N(n702), .A0(\ctrl/add_1_root_add_16_2/n48 ), .B0(
        \ctrl/add_1_root_add_16_2/n49 ), .Y(n405) );
  NAND2BX1 U864 ( .AN(\ctrl/add_1_root_add_16_2/n41 ), .B(
        \ctrl/add_1_root_add_16_2/n44 ), .Y(n406) );
  XOR2X1 U865 ( .A(n405), .B(n406), .Y(n407) );
  CLKNAND2X2 U866 ( .A(n554), .B(\ctrl/sub_0_root_add_0_root_sub_16/n31 ), .Y(
        n408) );
  XOR2X1 U867 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n32 ), .B(n408), .Y(n409) );
  CLKINVX1 U868 ( .A(n1043), .Y(n410) );
  AOI22XL U869 ( .A0(n1043), .A1(n407), .B0(n409), .B1(n410), .Y(D[25]) );
  AOI21X1 U870 ( .A0(n715), .A1(\normal/srl_15/n219 ), .B0(n504), .Y(n411) );
  OAI2B1X1 U871 ( .A1N(\normal/srl_15/n217 ), .A0(n715), .B0(n411), .Y(
        \normal/srl_15/n117 ) );
  AOI21X1 U872 ( .A0(n715), .A1(\normal/srl_15/n222 ), .B0(n504), .Y(n412) );
  OAI2B1X1 U873 ( .A1N(\normal/srl_15/n220 ), .A0(n715), .B0(n412), .Y(
        \normal/srl_15/n120 ) );
  AOI21X1 U874 ( .A0(n715), .A1(\normal/srl_15/n228 ), .B0(n504), .Y(n413) );
  OAI2B1X1 U875 ( .A1N(\normal/srl_15/n226 ), .A0(n715), .B0(n413), .Y(
        \normal/srl_15/n126 ) );
  AOI21X1 U876 ( .A0(n715), .A1(\normal/srl_15/n229 ), .B0(n504), .Y(n414) );
  OAI2B1X1 U877 ( .A1N(\normal/srl_15/n227 ), .A0(n715), .B0(n414), .Y(
        \normal/srl_15/n127 ) );
  AOI21X1 U878 ( .A0(n514), .A1(\normal/sll_15/n206 ), .B0(n504), .Y(n415) );
  OAI2B1X1 U879 ( .A1N(\normal/sll_15/n208 ), .A0(n514), .B0(n415), .Y(
        \normal/sll_15/n114 ) );
  CLKINVX1 U880 ( .A(\normal/sll_15/n1 ), .Y(n416) );
  CLKINVX1 U881 ( .A(n704), .Y(n417) );
  AOI22XL U882 ( .A0(n503), .A1(n416), .B0(\normal/sll_15/n49 ), .B1(n417), 
        .Y(n418) );
  OAI21X1 U883 ( .A0(n503), .A1(\normal/sll_15/n5 ), .B0(n418), .Y(n419) );
  OAI32XL U884 ( .A0(n419), .A1(\normal/sll_15/n51 ), .A2(\normal/sll_15/n50 ), 
        .B0(n417), .B1(n419), .Y(n997) );
  CLKINVX1 U885 ( .A(n503), .Y(n420) );
  AOI22XL U886 ( .A0(n503), .A1(\normal/srl_15/n36 ), .B0(\normal/srl_15/n35 ), 
        .B1(n420), .Y(n421) );
  AOI22XL U887 ( .A0(n503), .A1(\normal/sll_15/n34 ), .B0(\normal/sll_15/n35 ), 
        .B1(n420), .Y(n422) );
  MX2X1 U888 ( .A(n421), .B(n422), .S0(n999), .Y(norm_out[14]) );
  CLKINVX1 U889 ( .A(n503), .Y(n423) );
  AOI22XL U890 ( .A0(n503), .A1(\normal/srl_15/n38 ), .B0(\normal/srl_15/n37 ), 
        .B1(n423), .Y(n424) );
  AOI22XL U891 ( .A0(n503), .A1(\normal/sll_15/n36 ), .B0(\normal/sll_15/n37 ), 
        .B1(n423), .Y(n425) );
  MX2X1 U892 ( .A(n424), .B(n425), .S0(n999), .Y(norm_out[16]) );
  NOR3BX1 U893 ( .AN(\round/r298/n1 ), .B(\round/r298/n19 ), .C(
        \round/r298/n16 ), .Y(n426) );
  XOR2X1 U894 ( .A(norm_out[25]), .B(n426), .Y(\round/N30 ) );
  AOI222XL U895 ( .A0(n1026), .A1(norm_out[22]), .B0(n39), .B1(\round/N28 ), 
        .C0(n662), .C1(\round/N27 ), .Y(n427) );
  CLKINVX1 U896 ( .A(n427), .Y(D[19]) );
  CLKNAND2X2 U897 ( .A(n555), .B(\ctrl/sub_0_root_add_0_root_sub_16/n23 ), .Y(
        n428) );
  XOR2X1 U898 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n24 ), .B(n428), .Y(n429) );
  AOI21X1 U899 ( .A0(n702), .A1(\ctrl/add_1_root_add_16_2/n30 ), .B0(
        \ctrl/add_1_root_add_16_2/n31 ), .Y(n430) );
  CLKNAND2X2 U900 ( .A(n533), .B(\ctrl/add_1_root_add_16_2/n28 ), .Y(n431) );
  CLKNAND2X2 U901 ( .A(n430), .B(n431), .Y(n432) );
  OAI211XL U902 ( .A0(n431), .A1(n430), .B0(n432), .C0(n1043), .Y(n433) );
  OAI21X1 U903 ( .A0(n1043), .A1(n429), .B0(n433), .Y(D[27]) );
  AOI21X1 U904 ( .A0(n715), .A1(\normal/srl_15/n220 ), .B0(n504), .Y(n434) );
  OAI2B1X1 U905 ( .A1N(\normal/srl_15/n218 ), .A0(n715), .B0(n434), .Y(
        \normal/srl_15/n118 ) );
  AOI21X1 U906 ( .A0(n715), .A1(\normal/srl_15/n223 ), .B0(n504), .Y(n435) );
  OAI2B1X1 U907 ( .A1N(\normal/srl_15/n221 ), .A0(n715), .B0(n435), .Y(
        \normal/srl_15/n121 ) );
  AOI21X1 U908 ( .A0(n715), .A1(\normal/srl_15/n230 ), .B0(n504), .Y(n436) );
  OAI2B1X1 U909 ( .A1N(\normal/srl_15/n228 ), .A0(n715), .B0(n436), .Y(
        \normal/srl_15/n128 ) );
  AOI21X1 U910 ( .A0(n514), .A1(\normal/sll_15/n207 ), .B0(n504), .Y(n437) );
  OAI2B1X1 U911 ( .A1N(\normal/sll_15/n209 ), .A0(n514), .B0(n437), .Y(
        \normal/sll_15/n115 ) );
  NOR4BX1 U912 ( .AN(add_out[26]), .B(add_out[28]), .C(n956), .D(
        \normal/srl_15/A[27] ), .Y(n929) );
  OAI21X1 U913 ( .A0(\round/r298/n103 ), .A1(\round/r298/n104 ), .B0(
        norm_out[9]), .Y(n438) );
  OAI31X1 U914 ( .A0(\round/r298/n103 ), .A1(norm_out[9]), .A2(
        \round/r298/n104 ), .B0(n438), .Y(\round/N14 ) );
  CLKINVX1 U915 ( .A(n503), .Y(n439) );
  AOI22XL U916 ( .A0(n503), .A1(\normal/srl_15/n37 ), .B0(\normal/srl_15/n36 ), 
        .B1(n439), .Y(n440) );
  AOI22XL U917 ( .A0(n503), .A1(\normal/sll_15/n35 ), .B0(\normal/sll_15/n36 ), 
        .B1(n439), .Y(n441) );
  MX2X1 U918 ( .A(n440), .B(n441), .S0(n999), .Y(norm_out[15]) );
  CLKINVX1 U919 ( .A(n503), .Y(n442) );
  AOI22XL U920 ( .A0(n503), .A1(\normal/srl_15/n39 ), .B0(\normal/srl_15/n38 ), 
        .B1(n442), .Y(n443) );
  AOI22XL U921 ( .A0(n503), .A1(\normal/sll_15/n37 ), .B0(\normal/sll_15/n38 ), 
        .B1(n442), .Y(n444) );
  MX2X1 U922 ( .A(n443), .B(n444), .S0(n999), .Y(norm_out[17]) );
  NAND2BX1 U923 ( .AN(\round/r298/n31 ), .B(\round/r298/n1 ), .Y(n445) );
  XOR2X1 U924 ( .A(\round/r298/n28 ), .B(n445), .Y(\round/N27 ) );
  CLKINVX1 U925 ( .A(n503), .Y(n446) );
  AOI22XL U926 ( .A0(n503), .A1(\normal/srl_15/n47 ), .B0(\normal/srl_15/n46 ), 
        .B1(n446), .Y(n447) );
  AOI22XL U927 ( .A0(n503), .A1(\normal/sll_15/n45 ), .B0(\normal/sll_15/n46 ), 
        .B1(n446), .Y(n448) );
  MX2X1 U928 ( .A(n447), .B(n448), .S0(n999), .Y(norm_out[25]) );
  AOI222XL U929 ( .A0(n1026), .A1(norm_out[23]), .B0(n39), .B1(\round/N29 ), 
        .C0(n1025), .C1(\round/N28 ), .Y(n449) );
  CLKINVX1 U930 ( .A(n449), .Y(D[20]) );
  CLKNAND2X2 U931 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n36 ), .B(
        \ctrl/sub_0_root_add_0_root_sub_16/n14 ), .Y(n450) );
  XNOR2X1 U932 ( .A(n450), .B(\ctrl/sub_0_root_add_0_root_sub_16/n19 ), .Y(
        n451) );
  AOI21X1 U933 ( .A0(n702), .A1(\ctrl/add_1_root_add_16_2/n21 ), .B0(
        \ctrl/add_1_root_add_16_2/n22 ), .Y(n452) );
  CLKNAND2X2 U934 ( .A(\ctrl/add_1_root_add_16_2/n65 ), .B(
        \ctrl/add_1_root_add_16_2/n19 ), .Y(n453) );
  CLKNAND2X2 U935 ( .A(n452), .B(n453), .Y(n454) );
  OAI211XL U936 ( .A0(n453), .A1(n452), .B0(n454), .C0(n1043), .Y(n455) );
  OAI21X1 U937 ( .A0(n1043), .A1(n451), .B0(n455), .Y(D[28]) );
  AOI21X1 U938 ( .A0(n715), .A1(\normal/srl_15/n231 ), .B0(n504), .Y(n456) );
  OAI2B1X1 U939 ( .A1N(\normal/srl_15/n229 ), .A0(n715), .B0(n456), .Y(
        \normal/srl_15/n129 ) );
  AOI21X1 U940 ( .A0(n715), .A1(\normal/srl_15/n232 ), .B0(n504), .Y(n457) );
  OAI2B1X1 U941 ( .A1N(\normal/srl_15/n230 ), .A0(n715), .B0(n457), .Y(
        \normal/srl_15/n130 ) );
  AOI21X1 U942 ( .A0(n514), .A1(\normal/sll_15/n205 ), .B0(n504), .Y(n458) );
  OAI2B1X1 U943 ( .A1N(\normal/sll_15/n207 ), .A0(n514), .B0(n458), .Y(
        \normal/sll_15/n113 ) );
  AOI21X1 U944 ( .A0(n715), .A1(\normal/sll_15/n208 ), .B0(n504), .Y(n459) );
  OAI2B1X1 U945 ( .A1N(\normal/sll_15/n210 ), .A0(n715), .B0(n459), .Y(
        \normal/sll_15/n116 ) );
  CLKINVX1 U946 ( .A(n503), .Y(n460) );
  AOI22XL U947 ( .A0(n503), .A1(\normal/srl_15/n12 ), .B0(\normal/srl_15/n10 ), 
        .B1(n460), .Y(n461) );
  NOR4BX1 U948 ( .AN(\normal/srl_15/n11 ), .B(\normal/N14 ), .C(\normal/N15 ), 
        .D(n461), .Y(n462) );
  OAI21X1 U949 ( .A0(\normal/srl_15/n14 ), .A1(n503), .B0(\normal/srl_15/n15 ), 
        .Y(n463) );
  OAI21X1 U950 ( .A0(\normal/srl_15/n18 ), .A1(n460), .B0(\normal/srl_15/n17 ), 
        .Y(n464) );
  NOR3BX1 U951 ( .AN(\normal/srl_15/n16 ), .B(n463), .C(n464), .Y(n465) );
  NAND3XL U952 ( .A(n522), .B(n462), .C(n465), .Y(n990) );
  XOR2X1 U953 ( .A(norm_out[6]), .B(\round/r298/n112 ), .Y(\round/N11 ) );
  OAI21X1 U954 ( .A0(\round/r298/n95 ), .A1(\round/r298/n104 ), .B0(
        norm_out[10]), .Y(n466) );
  OAI31X1 U955 ( .A0(\round/r298/n95 ), .A1(norm_out[10]), .A2(
        \round/r298/n104 ), .B0(n466), .Y(\round/N15 ) );
  CLKINVX1 U956 ( .A(n503), .Y(n467) );
  AOI22XL U957 ( .A0(n503), .A1(\normal/srl_15/n34 ), .B0(\normal/srl_15/n33 ), 
        .B1(n467), .Y(n468) );
  AOI22XL U958 ( .A0(n503), .A1(\normal/sll_15/n32 ), .B0(\normal/sll_15/n33 ), 
        .B1(n467), .Y(n469) );
  MX2X1 U959 ( .A(n468), .B(n469), .S0(n999), .Y(norm_out[12]) );
  CLKINVX1 U960 ( .A(n503), .Y(n470) );
  AOI22XL U961 ( .A0(n503), .A1(\normal/srl_15/n40 ), .B0(\normal/srl_15/n39 ), 
        .B1(n470), .Y(n471) );
  AOI22XL U962 ( .A0(n503), .A1(\normal/sll_15/n38 ), .B0(\normal/sll_15/n39 ), 
        .B1(n470), .Y(n472) );
  MX2X1 U963 ( .A(n471), .B(n472), .S0(n999), .Y(norm_out[18]) );
  NOR3BX1 U964 ( .AN(\round/r298/n1 ), .B(\round/r298/n31 ), .C(
        \round/r298/n28 ), .Y(n473) );
  XOR2X1 U965 ( .A(norm_out[23]), .B(n473), .Y(\round/N28 ) );
  AOI21BX1 U966 ( .A0(n534), .A1(\ctrl/add_1_root_add_16_2/n60 ), .B0N(
        \ctrl/add_1_root_add_16_2/n57 ), .Y(\ctrl/add_1_root_add_16_2/n49 ) );
  AOI222XL U967 ( .A0(n1026), .A1(norm_out[24]), .B0(n39), .B1(\round/N30 ), 
        .C0(n1025), .C1(\round/N29 ), .Y(n474) );
  CLKINVX1 U968 ( .A(n474), .Y(D[21]) );
  XOR2X1 U969 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n12 ), .B(
        \ctrl/sub_0_root_add_0_root_sub_16/n10 ), .Y(n475) );
  CLKNAND2X2 U970 ( .A(\ctrl/add_1_root_add_16_2/n15 ), .B(n1034), .Y(n476) );
  OAI211XL U971 ( .A0(\ctrl/add_1_root_add_16_2/n15 ), .A1(n1034), .B0(n1043), 
        .C0(n476), .Y(n477) );
  OAI21X1 U972 ( .A0(n1043), .A1(n475), .B0(n477), .Y(D[29]) );
  AOI21X1 U973 ( .A0(n514), .A1(\normal/sll_15/n204 ), .B0(n504), .Y(n478) );
  OAI2B1X1 U974 ( .A1N(\normal/sll_15/n206 ), .A0(n514), .B0(n478), .Y(
        \normal/sll_15/n112 ) );
  AOI21X1 U975 ( .A0(n715), .A1(\normal/sll_15/n209 ), .B0(n504), .Y(n479) );
  OAI2B1X1 U976 ( .A1N(\normal/sll_15/n211 ), .A0(n715), .B0(n479), .Y(
        \normal/sll_15/n117 ) );
  AOI21X1 U977 ( .A0(n514), .A1(\normal/sll_15/n210 ), .B0(n504), .Y(n480) );
  OAI2B1X1 U978 ( .A1N(\normal/sll_15/n212 ), .A0(n514), .B0(n480), .Y(
        \normal/sll_15/n118 ) );
  NOR4X1 U979 ( .A(\normal/N8 ), .B(\normal/N9 ), .C(\normal/N10 ), .D(
        \normal/N11 ), .Y(n481) );
  NOR4X1 U980 ( .A(\normal/N4 ), .B(\normal/N5 ), .C(\normal/N6 ), .D(
        \normal/N7 ), .Y(n482) );
  NAND2BX1 U981 ( .AN(\normal/srl_15/n20 ), .B(n503), .Y(n483) );
  OAI211XL U982 ( .A0(n503), .A1(\normal/srl_15/n18 ), .B0(n483), .C0(
        \normal/srl_15/n19 ), .Y(n484) );
  NOR4X1 U983 ( .A(\normal/N22 ), .B(\normal/N23 ), .C(\normal/N3 ), .D(n484), 
        .Y(n485) );
  NAND3XL U984 ( .A(n481), .B(n482), .C(n485), .Y(n991) );
  XOR2X1 U985 ( .A(\round/r298/n116 ), .B(norm_out[5]), .Y(\round/N10 ) );
  CLKNAND2X2 U986 ( .A(\round/r298/n112 ), .B(norm_out[6]), .Y(n486) );
  XNOR2X1 U987 ( .A(n486), .B(norm_out[7]), .Y(\round/N12 ) );
  NOR3BX1 U988 ( .AN(norm_out[10]), .B(\round/r298/n95 ), .C(\round/r298/n104 ), .Y(n487) );
  XOR2X1 U989 ( .A(norm_out[11]), .B(n487), .Y(\round/N16 ) );
  CLKINVX1 U990 ( .A(n503), .Y(n488) );
  AOI22XL U991 ( .A0(n503), .A1(\normal/srl_15/n35 ), .B0(\normal/srl_15/n34 ), 
        .B1(n488), .Y(n489) );
  AOI22XL U992 ( .A0(n503), .A1(\normal/sll_15/n33 ), .B0(\normal/sll_15/n34 ), 
        .B1(n488), .Y(n490) );
  MX2X1 U993 ( .A(n489), .B(n490), .S0(n999), .Y(norm_out[13]) );
  CLKINVX1 U994 ( .A(n503), .Y(n491) );
  AOI22XL U995 ( .A0(n503), .A1(\normal/srl_15/n41 ), .B0(\normal/srl_15/n40 ), 
        .B1(n491), .Y(n492) );
  AOI22XL U996 ( .A0(n503), .A1(\normal/sll_15/n39 ), .B0(\normal/sll_15/n40 ), 
        .B1(n491), .Y(n493) );
  MX2X1 U997 ( .A(n492), .B(n493), .S0(n999), .Y(norm_out[19]) );
  OR2X1 U998 ( .A(n525), .B(\ctrl/add_1_root_add_16_2/n49 ), .Y(n494) );
  OAI211XL U999 ( .A0(\ctrl/add_1_root_add_16_2/n36 ), .A1(
        \ctrl/add_1_root_add_16_2/n44 ), .B0(\ctrl/add_1_root_add_16_2/n37 ), 
        .C0(n494), .Y(\ctrl/add_1_root_add_16_2/n31 ) );
  NOR3BX1 U1000 ( .AN(\round/r298/n1 ), .B(\round/r298/n9 ), .C(
        \round/r298/n19 ), .Y(n495) );
  XNOR2X1 U1001 ( .A(n556), .B(n495), .Y(n496) );
  AOI222XL U1002 ( .A0(n496), .A1(n39), .B0(n662), .B1(\round/N30 ), .C0(
        norm_out[25]), .C1(n1026), .Y(n497) );
  CLKINVX1 U1003 ( .A(n497), .Y(D[22]) );
  CLKNAND2X2 U1004 ( .A(\ctrl/add_1_root_add_16_2/n8 ), .B(
        \ctrl/add_1_root_add_16_2/n7 ), .Y(n498) );
  OAI211XL U1005 ( .A0(\ctrl/add_1_root_add_16_2/n8 ), .A1(
        \ctrl/add_1_root_add_16_2/n7 ), .B0(n1043), .C0(n498), .Y(n499) );
  XOR2X1 U1006 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n7 ), .B(
        \ctrl/sub_0_root_add_0_root_sub_16/A[7] ), .Y(n500) );
  OAI21X1 U1007 ( .A0(n1043), .A1(n500), .B0(n499), .Y(D[30]) );
  INVX2 U1008 ( .A(sig_B[0]), .Y(n678) );
  INVX2 U1009 ( .A(sig_A[2]), .Y(n669) );
  INVX2 U1010 ( .A(sig_A[5]), .Y(n668) );
  MXI2X8 U1011 ( .A(sig_P[49]), .B(\selc/N162 ), .S0(n775), .Y(n519) );
  MXI2X2 U1012 ( .A(\sub/r301/n17 ), .B(
        \expadd/add_0_root_sub_0_root_sub_8/n2 ), .S0(n516), .Y(
        \ctrl/add_1_root_add_16_2/A[0] ) );
  OAI21X1 U1013 ( .A0(n1002), .A1(n1001), .B0(n1000), .Y(n1003) );
  OAI21X1 U1014 ( .A0(n991), .A1(n990), .B0(n989), .Y(n1004) );
  MX2X1 U1015 ( .A(\normal/N45 ), .B(\normal/N91 ), .S0(n999), .Y(norm_out[23]) );
  MX2X1 U1016 ( .A(\normal/N33 ), .B(\normal/N79 ), .S0(n999), .Y(norm_out[11]) );
  MX2X1 U1017 ( .A(\normal/N27 ), .B(\normal/N73 ), .S0(n999), .Y(norm_out[5])
         );
  MX2X1 U1018 ( .A(\normal/N44 ), .B(\normal/N90 ), .S0(n999), .Y(norm_out[22]) );
  MX2X2 U1019 ( .A(\normal/N32 ), .B(\normal/N78 ), .S0(n999), .Y(norm_out[10]) );
  CLKBUFX24 U1020 ( .A(zero_cnt[0]), .Y(n503) );
  OAI21X2 U1021 ( .A0(n922), .A1(add_out[2]), .B0(n921), .Y(n967) );
  CLKINVX2 U1022 ( .A(n922), .Y(n906) );
  NAND2X2 U1023 ( .A(n864), .B(\normal/srl_15/A[1] ), .Y(n922) );
  INVX2 U1024 ( .A(n864), .Y(n881) );
  AOI21X1 U1025 ( .A0(n920), .A1(add_out[7]), .B0(n919), .Y(n921) );
  CLKNAND2X2 U1026 ( .A(\sigadd/N48 ), .B(n501), .Y(n788) );
  CLKNAND2X2 U1027 ( .A(\sigadd/N49 ), .B(n501), .Y(n830) );
  NAND2X2 U1028 ( .A(\sigadd/N19 ), .B(n501), .Y(n817) );
  CLKNAND2X2 U1029 ( .A(\sigadd/N50 ), .B(n501), .Y(n831) );
  NAND2X2 U1030 ( .A(\sigadd/N18 ), .B(n501), .Y(n818) );
  MX2X2 U1031 ( .A(\sigadd/sig[2] ), .B(\sigadd/N4 ), .S0(D[31]), .Y(
        add_out[2]) );
  CLKNAND2X2 U1032 ( .A(\sigadd/N46 ), .B(D[31]), .Y(n790) );
  MX2X2 U1033 ( .A(\sigadd/sig[4] ), .B(\sigadd/N6 ), .S0(D[31]), .Y(
        \normal/srl_15/A[4] ) );
  CLKNAND2X2 U1034 ( .A(\sigadd/N45 ), .B(D[31]), .Y(n791) );
  NAND2X2 U1035 ( .A(\sigadd/N31 ), .B(D[31]), .Y(n805) );
  CLKNAND2X2 U1036 ( .A(\sigadd/N47 ), .B(D[31]), .Y(n789) );
  INVX12 U1037 ( .A(n661), .Y(n501) );
  NAND2XL U1038 ( .A(\sigadd/N14 ), .B(\sigadd/sub_add_11_b0/B[49] ), .Y(n822)
         );
  INVX2 U1039 ( .A(\sigadd/add_9/n73 ), .Y(\sigadd/add_9/n71 ) );
  INVX2 U1040 ( .A(\sigadd/add_9/n65 ), .Y(\sigadd/add_9/n63 ) );
  MX2X1 U1041 ( .A(\align/N9 ), .B(sel_P[5]), .S0(n516), .Y(ali_P[5]) );
  MX2X1 U1042 ( .A(\align/N8 ), .B(sel_P[4]), .S0(n516), .Y(ali_P[4]) );
  MX2X1 U1043 ( .A(\align/N7 ), .B(sel_P[3]), .S0(n516), .Y(ali_P[3]) );
  CLKNAND2X2 U1044 ( .A(\selc/N147 ), .B(n502), .Y(n741) );
  CLKNAND2X2 U1045 ( .A(\selc/N146 ), .B(n502), .Y(n742) );
  CLKNAND2X2 U1046 ( .A(\selc/N145 ), .B(n502), .Y(n743) );
  NAND2X1 U1047 ( .A(\selc/N144 ), .B(n502), .Y(n744) );
  NAND2X1 U1048 ( .A(\selc/N143 ), .B(n502), .Y(n745) );
  NAND2XL U1049 ( .A(\selc/N142 ), .B(n502), .Y(n746) );
  NAND2XL U1050 ( .A(\selc/N141 ), .B(n502), .Y(n747) );
  NAND2XL U1051 ( .A(\selc/N140 ), .B(n502), .Y(n748) );
  CLKINVX1 U1052 ( .A(mux_out[7]), .Y(\ctrl/add_1_root_add_16_2/n7 ) );
  OA21XL U1053 ( .A0(\mul/mult_6/n1383 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n993 ), .Y(n607) );
  OAI21X4 U1054 ( .A0(\mul/mult_6/n623 ), .A1(\mul/mult_6/n575 ), .B0(
        \mul/mult_6/n576 ), .Y(\mul/mult_6/n1364 ) );
  OAI21X1 U1055 ( .A0(n678), .A1(\mul/mult_6/n76 ), .B0(n537), .Y(
        \mul/mult_6/n387 ) );
  BUFX3 U1056 ( .A(\mul/mult_6/n543 ), .Y(n700) );
  INVXL U1057 ( .A(\mul/mult_6/n683 ), .Y(\mul/mult_6/n726 ) );
  BUFX3 U1058 ( .A(\mul/mult_6/n547 ), .Y(n701) );
  INVX2 U1059 ( .A(sig_A[11]), .Y(n666) );
  INVX2 U1060 ( .A(sig_B[9]), .Y(n675) );
  INVX1 U1061 ( .A(sig_C[23]), .Y(\selc/r300/carry[24] ) );
  INVX2 U1062 ( .A(sig_B[21]), .Y(n670) );
  INVX6 U1063 ( .A(n1007), .Y(n1026) );
  INVXL U1064 ( .A(norm_out[17]), .Y(\round/r298/n56 ) );
  INVXL U1065 ( .A(norm_out[18]), .Y(\round/r298/n49 ) );
  INVXL U1066 ( .A(norm_out[12]), .Y(\round/r298/n83 ) );
  INVXL U1067 ( .A(norm_out[13]), .Y(\round/r298/n80 ) );
  BUFX12 U1068 ( .A(\normal/n30 ), .Y(n704) );
  CLKBUFX32 U1069 ( .A(zero_cnt[3]), .Y(n513) );
  NOR2X2 U1070 ( .A(\normal/srl_15/A[40] ), .B(add_out[39]), .Y(n948) );
  OAI21X2 U1071 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n588), .B0(n795), .Y(
        add_out[39]) );
  CLKNAND2X2 U1072 ( .A(\sigadd/N12 ), .B(n501), .Y(n824) );
  NAND2X1 U1073 ( .A(\sigadd/N13 ), .B(n501), .Y(n823) );
  OAI21X2 U1074 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n587), .B0(n793), .Y(
        \normal/srl_15/A[41] ) );
  OAI21X2 U1075 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n634), .B0(n822), .Y(
        \normal/srl_15/A[12] ) );
  BUFX10 U1076 ( .A(\sigadd/sub_add_11_b0/B[49] ), .Y(D[31]) );
  BUFX16 U1077 ( .A(\sigadd/n15 ), .Y(\sigadd/sub_add_11_b0/B[49] ) );
  INVX2 U1078 ( .A(\sigadd/add_9/n81 ), .Y(\sigadd/add_9/n79 ) );
  INVX2 U1079 ( .A(\sigadd/add_9/n89 ), .Y(\sigadd/add_9/n87 ) );
  INVX2 U1080 ( .A(\sigadd/add_9/n129 ), .Y(\sigadd/add_9/n127 ) );
  INVX2 U1081 ( .A(\sigadd/add_9/n121 ), .Y(\sigadd/add_9/n119 ) );
  INVX2 U1082 ( .A(\sigadd/add_9/n105 ), .Y(\sigadd/add_9/n103 ) );
  INVX2 U1083 ( .A(\sigadd/add_9/n97 ), .Y(\sigadd/add_9/n95 ) );
  INVX2 U1084 ( .A(\sigadd/add_9/n113 ), .Y(\sigadd/add_9/n111 ) );
  MX2X1 U1085 ( .A(\align/N12 ), .B(sel_P[8]), .S0(n516), .Y(ali_P[8]) );
  MX2X1 U1086 ( .A(\align/N11 ), .B(sel_P[7]), .S0(n516), .Y(ali_P[7]) );
  MX2X1 U1087 ( .A(\align/N10 ), .B(sel_P[6]), .S0(n516), .Y(ali_P[6]) );
  INVX2 U1088 ( .A(\mul/mult_6/n126 ), .Y(sig_P[49]) );
  INVX2 U1089 ( .A(sig_P[46]), .Y(\selc/r299/A[46] ) );
  NAND2XL U1090 ( .A(\selc/N139 ), .B(n502), .Y(n749) );
  NAND2XL U1091 ( .A(\selc/N138 ), .B(n502), .Y(n750) );
  NAND2XL U1092 ( .A(\selc/N137 ), .B(n502), .Y(n751) );
  NAND2XL U1093 ( .A(\selc/N136 ), .B(n502), .Y(n752) );
  NAND2XL U1094 ( .A(\selc/N135 ), .B(n502), .Y(n753) );
  NAND2XL U1095 ( .A(\selc/N134 ), .B(n502), .Y(n754) );
  NAND2XL U1096 ( .A(\selc/N133 ), .B(n502), .Y(n755) );
  NAND2XL U1097 ( .A(\selc/N132 ), .B(n502), .Y(n756) );
  CLKNAND2X2 U1098 ( .A(exp_P[7]), .B(n1027), .Y(n782) );
  CLKNAND2X2 U1099 ( .A(n778), .B(n777), .Y(n784) );
  OA21XL U1100 ( .A0(\mul/mult_6/n1382 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n992 ), .Y(n628) );
  BUFX5 U1101 ( .A(\mul/mult_6/n42 ), .Y(n687) );
  BUFX5 U1102 ( .A(\mul/mult_6/n22 ), .Y(n683) );
  BUFX3 U1103 ( .A(\mul/mult_6/n539 ), .Y(n699) );
  BUFX5 U1104 ( .A(\mul/mult_6/n32 ), .Y(n685) );
  INVX2 U1105 ( .A(sig_B[7]), .Y(n676) );
  INVX2 U1106 ( .A(sig_A[8]), .Y(n667) );
  INVXL U1107 ( .A(norm_out[19]), .Y(\round/r298/n44 ) );
  INVXL U1108 ( .A(norm_out[21]), .Y(\round/r298/n35 ) );
  BUFX12 U1109 ( .A(\normal/n30 ), .Y(n512) );
  BUFX16 U1110 ( .A(zero_cnt[4]), .Y(n703) );
  NOR2X2 U1111 ( .A(n944), .B(add_out[45]), .Y(n833) );
  NOR2X2 U1112 ( .A(add_out[16]), .B(add_out[17]), .Y(n873) );
  OAI21X2 U1113 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n633), .B0(n820), .Y(
        add_out[14]) );
  INVX2 U1114 ( .A(\normal/srl_15/A[41] ), .Y(n834) );
  CLKNAND2X2 U1115 ( .A(\sigadd/N10 ), .B(n501), .Y(n826) );
  NAND2X1 U1116 ( .A(\sigadd/N11 ), .B(n501), .Y(n825) );
  CLKNAND2X2 U1117 ( .A(\sigadd/N15 ), .B(n501), .Y(n821) );
  NAND2XL U1118 ( .A(\sigadd/N8 ), .B(n501), .Y(n828) );
  OAI21X4 U1119 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n601), .B0(n804), .Y(
        add_out[30]) );
  OAI21X4 U1120 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n613), .B0(n805), .Y(
        \normal/srl_15/A[29] ) );
  OAI21X2 U1121 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n589), .B0(n797), .Y(
        add_out[37]) );
  OAI21X2 U1122 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n559), .B0(n790), .Y(
        \normal/srl_15/A[44] ) );
  OAI21X2 U1123 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n567), .B0(n791), .Y(
        add_out[43]) );
  XNOR2X1 U1124 ( .A(\sigadd/add_9/n61 ), .B(\sigadd/add_9/n3 ), .Y(n568) );
  XNOR2X1 U1125 ( .A(\sigadd/add_9/n85 ), .B(\sigadd/add_9/n9 ), .Y(n587) );
  XOR2X1 U1126 ( .A(\sigadd/add_9/n90 ), .B(\sigadd/add_9/n10 ), .Y(n581) );
  XNOR2X1 U1127 ( .A(\sigadd/add_9/n93 ), .B(\sigadd/add_9/n11 ), .Y(n588) );
  XOR2X1 U1128 ( .A(\sigadd/add_9/n98 ), .B(\sigadd/add_9/n12 ), .Y(n582) );
  XNOR2X1 U1129 ( .A(\sigadd/add_9/n101 ), .B(\sigadd/add_9/n13 ), .Y(n589) );
  XOR2X1 U1130 ( .A(\sigadd/add_9/n106 ), .B(\sigadd/add_9/n14 ), .Y(n583) );
  XNOR2X1 U1131 ( .A(\sigadd/add_9/n109 ), .B(\sigadd/add_9/n15 ), .Y(n590) );
  INVX2 U1132 ( .A(\sigadd/add_9/n57 ), .Y(\sigadd/add_9/n55 ) );
  MX2X1 U1133 ( .A(\align/N15 ), .B(sel_P[11]), .S0(n516), .Y(ali_P[11]) );
  MX2X1 U1134 ( .A(\align/N14 ), .B(sel_P[10]), .S0(n516), .Y(ali_P[10]) );
  MX2X1 U1135 ( .A(\align/N13 ), .B(sel_P[9]), .S0(n516), .Y(ali_P[9]) );
  MX2X1 U1136 ( .A(\align/N17 ), .B(sel_P[13]), .S0(n516), .Y(ali_P[13]) );
  MX2X1 U1137 ( .A(\align/N16 ), .B(sel_P[12]), .S0(n1030), .Y(ali_P[12]) );
  MXI2X1 U1138 ( .A(\align/sra_10/n191 ), .B(\align/sra_10/n195 ), .S0(n505), 
        .Y(\align/sra_10/n141 ) );
  OAI21X1 U1139 ( .A0(n502), .A1(\selc/r299/A[47] ), .B0(n728), .Y(sel_P[47])
         );
  OAI21X1 U1140 ( .A0(n502), .A1(\selc/r299/A[46] ), .B0(n729), .Y(sel_P[46])
         );
  ADDFX2 U1141 ( .A(\mul/mult_6/n180 ), .B(n670), .CI(\mul/mult_6/n128 ), .CO(
        \mul/mult_6/n127 ), .S(sig_P[47]) );
  ADDFX2 U1142 ( .A(\mul/mult_6/n253 ), .B(\mul/mult_6/n261 ), .CI(
        \mul/mult_6/n142 ), .CO(\mul/mult_6/n141 ), .S(sig_P[33]) );
  ADDFX2 U1143 ( .A(\mul/mult_6/n271 ), .B(\mul/mult_6/n280 ), .CI(
        \mul/mult_6/n144 ), .CO(\mul/mult_6/n143 ), .S(sig_P[31]) );
  ADDFX2 U1144 ( .A(\mul/mult_6/n346 ), .B(\mul/mult_6/n356 ), .CI(
        \mul/mult_6/n151 ), .CO(\mul/mult_6/n150 ), .S(sig_P[24]) );
  ADDFX2 U1145 ( .A(\mul/mult_6/n368 ), .B(\mul/mult_6/n378 ), .CI(
        \mul/mult_6/n153 ), .CO(\mul/mult_6/n152 ), .S(sig_P[22]) );
  NAND2XL U1146 ( .A(\selc/N131 ), .B(n724), .Y(n757) );
  NAND2XL U1147 ( .A(\selc/N130 ), .B(n502), .Y(n758) );
  NAND2XL U1148 ( .A(\selc/N129 ), .B(n502), .Y(n759) );
  NAND2XL U1149 ( .A(\selc/N127 ), .B(n502), .Y(n761) );
  OA21XL U1150 ( .A0(\mul/mult_6/n1375 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n985 ), .Y(n638) );
  OA21XL U1151 ( .A0(\mul/mult_6/n1380 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n990 ), .Y(n624) );
  OA21XL U1152 ( .A0(n542), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n988 ), .Y(
        n626) );
  OA21XL U1153 ( .A0(n572), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n986 ), .Y(
        n642) );
  OA21XL U1154 ( .A0(n543), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n989 ), .Y(
        n627) );
  OA21XL U1155 ( .A0(n544), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n991 ), .Y(
        n625) );
  OAI21X1 U1156 ( .A0(exp_P[3]), .A1(n1049), .B0(n726), .Y(n1052) );
  OA21XL U1157 ( .A0(n545), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n994 ), .Y(
        n605) );
  INVX2 U1158 ( .A(\mul/mult_6/n623 ), .Y(\mul/mult_6/n622 ) );
  OAI21XL U1159 ( .A0(exp_P[0]), .A1(\sub/r301/n17 ), .B0(n1044), .Y(n776) );
  BUFX5 U1160 ( .A(\mul/mult_6/n72 ), .Y(n695) );
  BUFX3 U1161 ( .A(\mul/mult_6/n54 ), .Y(n690) );
  OR2X2 U1162 ( .A(exp_P[0]), .B(\sub/r301/n17 ), .Y(n659) );
  BUFX5 U1163 ( .A(\mul/mult_6/n52 ), .Y(n689) );
  BUFX3 U1164 ( .A(\mul/mult_6/n535 ), .Y(n698) );
  NOR2BX4 U1165 ( .AN(\mul/mult_6/n1436 ), .B(\mul/mult_6/n1444 ), .Y(
        \mul/mult_6/n74 ) );
  NOR2X2 U1166 ( .A(\mul/mult_6/n1436 ), .B(\mul/mult_6/n1452 ), .Y(
        \mul/mult_6/n72 ) );
  BUFX18 U1167 ( .A(n724), .Y(n502) );
  BUFX3 U1168 ( .A(\mul/mult_6/n64 ), .Y(n693) );
  INVX2 U1169 ( .A(sig_B[18]), .Y(n671) );
  INVX2 U1170 ( .A(sig_A[20]), .Y(n663) );
  INVX2 U1171 ( .A(sig_B[15]), .Y(n672) );
  INVX2 U1172 ( .A(sig_A[14]), .Y(n665) );
  INVX2 U1173 ( .A(sig_A[22]), .Y(\mul/mult_6/n1452 ) );
  XOR2X1 U1174 ( .A(sign_B), .B(sign_A), .Y(n775) );
  NAND2X1 U1175 ( .A(n39), .B(\round/N9 ), .Y(n1005) );
  INVX2 U1176 ( .A(\round/r298/n105 ), .Y(\round/r298/n104 ) );
  NAND2X4 U1177 ( .A(n1004), .B(n1003), .Y(n1007) );
  AND2X2 U1178 ( .A(\round/r298/n5 ), .B(\round/r298/n18 ), .Y(n563) );
  INVXL U1179 ( .A(\round/r298/n76 ), .Y(\round/r298/n75 ) );
  CLKINVX2 U1180 ( .A(\ctrl/add_1_root_add_16_2/n23 ), .Y(
        \ctrl/add_1_root_add_16_2/n21 ) );
  AND2X4 U1181 ( .A(n988), .B(n987), .Y(n522) );
  INVXL U1182 ( .A(norm_out[15]), .Y(\round/r298/n68 ) );
  OR3X6 U1183 ( .A(n967), .B(n937), .C(n936), .Y(\normal/n30 ) );
  INVX2 U1184 ( .A(n967), .Y(n986) );
  BUFX20 U1185 ( .A(zero_cnt[1]), .Y(n514) );
  NOR2X6 U1186 ( .A(n903), .B(n850), .Y(n864) );
  OAI21X1 U1187 ( .A0(n964), .A1(n918), .B0(n917), .Y(n919) );
  BUFX8 U1188 ( .A(zero_cnt[4]), .Y(n714) );
  NOR2X2 U1189 ( .A(n853), .B(n852), .Y(n982) );
  NAND2X6 U1190 ( .A(n875), .B(n844), .Y(n980) );
  NAND2X6 U1191 ( .A(n909), .B(n834), .Y(n949) );
  INVX2 U1192 ( .A(add_out[19]), .Y(n979) );
  NOR3X4 U1193 ( .A(add_out[46]), .B(add_out[47]), .C(add_out[49]), .Y(n832)
         );
  OAI21X2 U1194 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n646), .B0(n823), .Y(
        \normal/srl_15/A[11] ) );
  OAI21X2 U1195 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n612), .B0(n803), .Y(
        add_out[31]) );
  OAI21X2 U1196 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n600), .B0(n802), .Y(
        \normal/srl_15/A[32] ) );
  MX2X2 U1197 ( .A(\sigadd/sig[3] ), .B(\sigadd/N5 ), .S0(D[31]), .Y(
        add_out[3]) );
  MX2X2 U1198 ( .A(\sigadd/sig[1] ), .B(\sigadd/N3 ), .S0(D[31]), .Y(
        \normal/srl_15/A[1] ) );
  NAND2X1 U1199 ( .A(\sigadd/N17 ), .B(\sigadd/sub_add_11_b0/B[49] ), .Y(n819)
         );
  NAND2XL U1200 ( .A(\sigadd/N9 ), .B(\sigadd/sub_add_11_b0/B[49] ), .Y(n827)
         );
  MXI2X2 U1201 ( .A(n656), .B(n829), .S0(\sigadd/sub_add_11_b0/B[49] ), .Y(
        add_out[5]) );
  XOR2X2 U1202 ( .A(\sigadd/add_9/n53 ), .B(\sigadd/add_9/n1 ), .Y(
        \sigadd/n15 ) );
  XOR2X1 U1203 ( .A(\sigadd/add_9/n58 ), .B(\sigadd/add_9/n2 ), .Y(n560) );
  XOR2X1 U1204 ( .A(\sigadd/add_9/n66 ), .B(\sigadd/add_9/n4 ), .Y(n558) );
  XNOR2X1 U1205 ( .A(\sigadd/add_9/n69 ), .B(\sigadd/add_9/n5 ), .Y(n566) );
  XOR2X1 U1206 ( .A(\sigadd/add_9/n74 ), .B(\sigadd/add_9/n6 ), .Y(n559) );
  XOR2X1 U1207 ( .A(\sigadd/add_9/n82 ), .B(\sigadd/add_9/n8 ), .Y(n580) );
  MX2X1 U1208 ( .A(\align/N23 ), .B(sel_P[19]), .S0(n516), .Y(ali_P[19]) );
  MX2X1 U1209 ( .A(\align/N25 ), .B(sel_P[21]), .S0(n516), .Y(ali_P[21]) );
  MX2X1 U1210 ( .A(\align/N22 ), .B(sel_P[18]), .S0(n516), .Y(ali_P[18]) );
  MX2X1 U1211 ( .A(\align/N21 ), .B(sel_P[17]), .S0(n516), .Y(ali_P[17]) );
  MX2X1 U1212 ( .A(\align/N24 ), .B(sel_P[20]), .S0(n516), .Y(ali_P[20]) );
  MX2X1 U1213 ( .A(\align/N20 ), .B(sel_P[16]), .S0(n516), .Y(ali_P[16]) );
  MX2X1 U1214 ( .A(\align/N19 ), .B(sel_P[15]), .S0(n516), .Y(ali_P[15]) );
  MX2X1 U1215 ( .A(\align/N18 ), .B(sel_P[14]), .S0(n516), .Y(ali_P[14]) );
  MXI2X1 U1216 ( .A(\align/sra_10/n185 ), .B(\align/sra_10/n189 ), .S0(n505), 
        .Y(\align/sra_10/n135 ) );
  INVX20 U1217 ( .A(n519), .Y(n706) );
  OAI21X1 U1218 ( .A0(n502), .A1(\selc/r299/A[45] ), .B0(n730), .Y(sel_P[45])
         );
  XOR2X2 U1219 ( .A(\mul/mult_6/n127 ), .B(sig_B[21]), .Y(n557) );
  OAI21X1 U1220 ( .A0(n502), .A1(\selc/r299/A[44] ), .B0(n731), .Y(sel_P[44])
         );
  OAI21X1 U1221 ( .A0(n502), .A1(\selc/r299/A[43] ), .B0(n732), .Y(sel_P[43])
         );
  OAI21X1 U1222 ( .A0(n502), .A1(\selc/r299/A[42] ), .B0(n733), .Y(sel_P[42])
         );
  OAI21X1 U1223 ( .A0(n502), .A1(\selc/r299/A[41] ), .B0(n734), .Y(sel_P[41])
         );
  OAI21X1 U1224 ( .A0(n502), .A1(\selc/r299/A[40] ), .B0(n735), .Y(sel_P[40])
         );
  ADDFX2 U1225 ( .A(\mul/mult_6/n190 ), .B(\mul/mult_6/n188 ), .CI(
        \mul/mult_6/n131 ), .CO(\mul/mult_6/n130 ), .S(sig_P[44]) );
  OAI21X1 U1226 ( .A0(n502), .A1(\selc/r299/A[39] ), .B0(n736), .Y(sel_P[39])
         );
  OAI21X1 U1227 ( .A0(n502), .A1(\selc/r299/A[38] ), .B0(n737), .Y(sel_P[38])
         );
  OAI21X1 U1228 ( .A0(n502), .A1(\selc/r299/A[37] ), .B0(n738), .Y(sel_P[37])
         );
  OAI21X1 U1229 ( .A0(n502), .A1(\selc/r299/A[36] ), .B0(n739), .Y(sel_P[36])
         );
  OAI21X1 U1230 ( .A0(n502), .A1(\selc/r299/A[35] ), .B0(n740), .Y(sel_P[35])
         );
  NAND2XL U1231 ( .A(\selc/N128 ), .B(n502), .Y(n760) );
  NAND2XL U1232 ( .A(\selc/N125 ), .B(n502), .Y(n763) );
  INVX2 U1233 ( .A(\align/sra_11/n667 ), .Y(n716) );
  MX2X1 U1234 ( .A(\sub/N19 ), .B(\sub/N10 ), .S0(n516), .Y(sub_out[5]) );
  OA21XL U1235 ( .A0(\mul/mult_6/n1367 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n977 ), .Y(n655) );
  OA21XL U1236 ( .A0(\mul/mult_6/n1369 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n979 ), .Y(n651) );
  OA21XL U1237 ( .A0(\mul/mult_6/n1373 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n983 ), .Y(n641) );
  OA21XL U1238 ( .A0(\mul/mult_6/n1377 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n987 ), .Y(n629) );
  OA21XL U1239 ( .A0(\mul/mult_6/n1366 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n976 ), .Y(n654) );
  OA21XL U1240 ( .A0(n571), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n984 ), .Y(
        n637) );
  OA21XL U1241 ( .A0(n591), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n978 ), .Y(
        n650) );
  OA21XL U1242 ( .A0(n570), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n982 ), .Y(
        n639) );
  OA21XL U1243 ( .A0(n569), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n980 ), .Y(
        n652) );
  ADDHX1 U1244 ( .A(sig_A[5]), .B(\mul/mult_6/n919 ), .CO(\mul/mult_6/n494 ), 
        .S(\mul/mult_6/n495 ) );
  OAI21X1 U1245 ( .A0(n678), .A1(\mul/mult_6/n18 ), .B0(n565), .Y(
        \mul/mult_6/n1284 ) );
  NAND2X2 U1246 ( .A(n681), .B(sig_B[0]), .Y(n565) );
  NOR2X2 U1247 ( .A(n1057), .B(n1058), .Y(n1059) );
  NOR2X2 U1248 ( .A(n1054), .B(n1055), .Y(n1056) );
  NOR2X6 U1249 ( .A(n521), .B(n1026), .Y(n1025) );
  NOR2X6 U1250 ( .A(n521), .B(n1026), .Y(n662) );
  MXI2X1 U1251 ( .A(\normal/N48 ), .B(\normal/N94 ), .S0(n999), .Y(n556) );
  OR3X2 U1252 ( .A(n937), .B(n906), .C(n905), .Y(zero_cnt[3]) );
  AOI211X2 U1253 ( .A0(n983), .A1(add_out[13]), .B0(n982), .C0(n981), .Y(n984)
         );
  INVX1 U1254 ( .A(n968), .Y(n983) );
  INVXL U1255 ( .A(n931), .Y(n932) );
  OAI31X1 U1256 ( .A0(n898), .A1(add_out[38]), .A2(n897), .B0(n896), .Y(n899)
         );
  OR3X1 U1257 ( .A(n913), .B(n869), .C(\normal/srl_15/A[25] ), .Y(n870) );
  INVX4 U1258 ( .A(add_out[48]), .Y(n972) );
  OAI21X2 U1259 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n649), .B0(n828), .Y(
        \normal/srl_15/A[6] ) );
  OAI21X4 U1260 ( .A0(n501), .A1(n615), .B0(n809), .Y(\normal/srl_15/A[25] )
         );
  NOR2X2 U1261 ( .A(add_out[38]), .B(add_out[37]), .Y(n835) );
  INVX2 U1262 ( .A(\normal/srl_15/A[12] ), .Y(n938) );
  OAI21X4 U1263 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n648), .B0(n827), .Y(
        add_out[7]) );
  INVX2 U1264 ( .A(\sigadd/add_9/n193 ), .Y(\sigadd/add_9/n191 ) );
  INVX2 U1265 ( .A(\sigadd/add_9/n201 ), .Y(\sigadd/add_9/n199 ) );
  INVX2 U1266 ( .A(\sigadd/add_9/n185 ), .Y(\sigadd/add_9/n183 ) );
  MX2X1 U1267 ( .A(\align/N29 ), .B(sel_P[25]), .S0(n516), .Y(ali_P[25]) );
  MX2X1 U1268 ( .A(\align/N27 ), .B(sel_P[23]), .S0(n516), .Y(ali_P[23]) );
  MX2X1 U1269 ( .A(\align/N26 ), .B(sel_P[22]), .S0(n516), .Y(ali_P[22]) );
  MXI2X1 U1270 ( .A(\align/sra_10/n193 ), .B(\align/sra_10/n197 ), .S0(n505), 
        .Y(\align/sra_10/n143 ) );
  MXI2X1 U1271 ( .A(\align/sra_10/n197 ), .B(n508), .S0(n505), .Y(
        \align/sra_10/n147 ) );
  MXI2X1 U1272 ( .A(\align/sra_10/n196 ), .B(\align/sra_10/n200 ), .S0(n505), 
        .Y(\align/sra_10/n146 ) );
  MXI2X1 U1273 ( .A(\align/sra_10/n195 ), .B(\align/sra_10/n199 ), .S0(n505), 
        .Y(\align/sra_10/n145 ) );
  MXI2X1 U1274 ( .A(\align/sra_10/n194 ), .B(\align/sra_10/n198 ), .S0(n505), 
        .Y(\align/sra_10/n144 ) );
  MXI2X1 U1275 ( .A(\align/sra_10/n189 ), .B(\align/sra_10/n193 ), .S0(n505), 
        .Y(\align/sra_10/n139 ) );
  OR2XL U1276 ( .A(n706), .B(\two_en[1] ), .Y(n539) );
  ADDHX2 U1277 ( .A(\selc/r299/n2 ), .B(n557), .CO(\selc/r299/n1 ), .S(
        \selc/N161 ) );
  ADDHX2 U1278 ( .A(\selc/r299/n3 ), .B(\selc/r299/A[47] ), .CO(\selc/r299/n2 ), .S(\selc/N160 ) );
  INVX2 U1279 ( .A(sig_P[45]), .Y(\selc/r299/A[45] ) );
  INVX2 U1280 ( .A(sig_P[44]), .Y(\selc/r299/A[44] ) );
  INVX2 U1281 ( .A(sig_P[43]), .Y(\selc/r299/A[43] ) );
  INVX2 U1282 ( .A(sig_P[42]), .Y(\selc/r299/A[42] ) );
  ADDFX2 U1283 ( .A(\mul/mult_6/n458 ), .B(\mul/mult_6/n464 ), .CI(
        \mul/mult_6/n163 ), .CO(\mul/mult_6/n162 ), .S(sig_P[12]) );
  BUFX12 U1284 ( .A(\align/sra_10/n254 ), .Y(n509) );
  INVX2 U1285 ( .A(\ctrl/add_1_root_add_16_2/A[2] ), .Y(n1040) );
  BUFX12 U1286 ( .A(sub_out[2]), .Y(n511) );
  CMPR42X1 U1287 ( .A(\mul/mult_6/n385 ), .B(\mul/mult_6/n391 ), .C(
        \mul/mult_6/n392 ), .D(\mul/mult_6/n382 ), .ICI(\mul/mult_6/n388 ), 
        .S(\mul/mult_6/n379 ), .ICO(\mul/mult_6/n377 ), .CO(\mul/mult_6/n378 )
         );
  CMPR42X1 U1288 ( .A(\mul/mult_6/n362 ), .B(\mul/mult_6/n352 ), .C(
        \mul/mult_6/n359 ), .D(\mul/mult_6/n349 ), .ICI(\mul/mult_6/n355 ), 
        .S(\mul/mult_6/n346 ), .ICO(\mul/mult_6/n344 ), .CO(\mul/mult_6/n345 )
         );
  CMPR42X1 U1289 ( .A(\mul/mult_6/n928 ), .B(\mul/mult_6/n904 ), .C(
        \mul/mult_6/n422 ), .D(\mul/mult_6/n413 ), .ICI(\mul/mult_6/n418 ), 
        .S(\mul/mult_6/n410 ), .ICO(\mul/mult_6/n408 ), .CO(\mul/mult_6/n409 )
         );
  OA21XL U1290 ( .A0(\mul/mult_6/n1371 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n981 ), .Y(n643) );
  OA21XL U1291 ( .A0(\mul/mult_6/n1365 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n975 ), .Y(n658) );
  OA21XL U1292 ( .A0(\mul/mult_6/n1363 ), .A1(\mul/mult_6/n76 ), .B0(n697), 
        .Y(n540) );
  OA21XL U1293 ( .A0(\mul/mult_6/n1364 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n974 ), .Y(n541) );
  NAND2X2 U1294 ( .A(n683), .B(sig_B[0]), .Y(n532) );
  INVX2 U1295 ( .A(\mul/mult_6/n699 ), .Y(\mul/mult_6/n698 ) );
  BUFX10 U1296 ( .A(\mul/mult_6/n2 ), .Y(n679) );
  INVX2 U1297 ( .A(\mul/mult_6/n707 ), .Y(\mul/mult_6/n708 ) );
  MX2X1 U1298 ( .A(\ctrl/N30 ), .B(\ctrl/N14 ), .S0(n1043), .Y(D[26]) );
  MX2X1 U1299 ( .A(\ctrl/N28 ), .B(\ctrl/N12 ), .S0(n1043), .Y(D[24]) );
  AOI21X2 U1300 ( .A0(n1040), .A1(n1041), .B0(n1039), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/A[2] ) );
  AND2X6 U1301 ( .A(n39), .B(\ctrl/add_1_root_add_16_2/A[0] ), .Y(n1042) );
  NOR4X2 U1302 ( .A(\normal/N58 ), .B(\normal/N59 ), .C(\normal/N60 ), .D(
        \normal/N61 ), .Y(n993) );
  INVX2 U1303 ( .A(norm_out[4]), .Y(\round/r298/n117 ) );
  NOR4X2 U1304 ( .A(\normal/N62 ), .B(\normal/N63 ), .C(\normal/N64 ), .D(
        \normal/N65 ), .Y(n992) );
  MXI2X1 U1305 ( .A(\normal/sll_15/n176 ), .B(\normal/sll_15/n144 ), .S0(n504), 
        .Y(\normal/sll_15/n129 ) );
  CLKBUFX32 U1306 ( .A(\normal/n29 ), .Y(n504) );
  BUFX20 U1307 ( .A(zero_cnt[1]), .Y(n715) );
  OAI211X2 U1308 ( .A0(n866), .A1(n881), .B0(n865), .C0(n922), .Y(\normal/n29 ) );
  OAI211X2 U1309 ( .A0(n903), .A1(n857), .B0(n856), .C0(n855), .Y(n966) );
  NOR2X4 U1310 ( .A(n964), .B(\normal/srl_15/A[8] ), .Y(n920) );
  OAI21X1 U1311 ( .A0(add_out[16]), .A1(add_out[18]), .B0(n932), .Y(n933) );
  INVXL U1312 ( .A(n940), .Y(n916) );
  NOR2X2 U1313 ( .A(n874), .B(\normal/srl_15/A[27] ), .Y(n841) );
  NOR2X2 U1314 ( .A(n943), .B(add_out[33]), .Y(n838) );
  INVX2 U1315 ( .A(\normal/srl_15/A[22] ), .Y(n889) );
  INVX2 U1316 ( .A(add_out[14]), .Y(n846) );
  INVX2 U1317 ( .A(\normal/srl_15/A[25] ), .Y(n842) );
  INVX2 U1318 ( .A(add_out[18]), .Y(n845) );
  NOR2X2 U1319 ( .A(add_out[24]), .B(add_out[23]), .Y(n869) );
  NOR2X2 U1320 ( .A(add_out[20]), .B(\normal/srl_15/A[21] ), .Y(n844) );
  INVX2 U1321 ( .A(\normal/srl_15/A[10] ), .Y(n848) );
  OAI21X4 U1322 ( .A0(n501), .A1(n604), .B0(n810), .Y(add_out[24]) );
  OAI21X4 U1323 ( .A0(n501), .A1(n621), .B0(n814), .Y(add_out[20]) );
  OAI21X4 U1324 ( .A0(n501), .A1(n630), .B0(n813), .Y(\normal/srl_15/A[21] )
         );
  OAI21X4 U1325 ( .A0(n501), .A1(n622), .B0(n816), .Y(add_out[18]) );
  OAI21X4 U1326 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n644), .B0(n819), .Y(
        add_out[15]) );
  INVX2 U1327 ( .A(add_out[5]), .Y(n894) );
  ADDHX2 U1328 ( .A(n612), .B(\sigadd/sub_add_11_b0/n19 ), .CO(
        \sigadd/sub_add_11_b0/n18 ), .S(\sigadd/N33 ) );
  ADDHX2 U1329 ( .A(n601), .B(\sigadd/sub_add_11_b0/n20 ), .CO(
        \sigadd/sub_add_11_b0/n19 ), .S(\sigadd/N32 ) );
  ADDHX2 U1330 ( .A(n614), .B(\sigadd/sub_add_11_b0/n23 ), .CO(
        \sigadd/sub_add_11_b0/n22 ), .S(\sigadd/N29 ) );
  ADDHX2 U1331 ( .A(n603), .B(\sigadd/sub_add_11_b0/n24 ), .CO(
        \sigadd/sub_add_11_b0/n23 ), .S(\sigadd/N28 ) );
  INVX2 U1332 ( .A(\sigadd/add_9/n161 ), .Y(\sigadd/add_9/n159 ) );
  INVX2 U1333 ( .A(\sigadd/add_9/n145 ), .Y(\sigadd/add_9/n143 ) );
  INVX2 U1334 ( .A(\sigadd/add_9/n153 ), .Y(\sigadd/add_9/n151 ) );
  INVX2 U1335 ( .A(\sigadd/add_9/n169 ), .Y(\sigadd/add_9/n167 ) );
  INVX2 U1336 ( .A(\sigadd/add_9/n177 ), .Y(\sigadd/add_9/n175 ) );
  INVX2 U1337 ( .A(\sigadd/add_9/n137 ), .Y(\sigadd/add_9/n135 ) );
  OR2XL U1338 ( .A(ali_P[0]), .B(ali_C[0]), .Y(n561) );
  MX2X1 U1339 ( .A(\align/N30 ), .B(sel_P[26]), .S0(n516), .Y(ali_P[26]) );
  MX2X1 U1340 ( .A(\align/N28 ), .B(sel_P[24]), .S0(n516), .Y(ali_P[24]) );
  MX2X1 U1341 ( .A(\align/N39 ), .B(sel_P[35]), .S0(n1030), .Y(ali_P[35]) );
  MX2X1 U1342 ( .A(\align/N47 ), .B(sel_P[43]), .S0(n516), .Y(ali_P[43]) );
  MX2X1 U1343 ( .A(\align/N38 ), .B(sel_P[34]), .S0(n1030), .Y(ali_P[34]) );
  MX2X1 U1344 ( .A(\align/N36 ), .B(sel_P[32]), .S0(n1030), .Y(ali_P[32]) );
  MX2X1 U1345 ( .A(\align/N52 ), .B(sel_P[48]), .S0(n516), .Y(ali_P[48]) );
  MX2X1 U1346 ( .A(\align/N37 ), .B(sel_P[33]), .S0(n1030), .Y(ali_P[33]) );
  MX2X1 U1347 ( .A(\align/N4 ), .B(sig_P[0]), .S0(n516), .Y(ali_P[0]) );
  MX2X1 U1348 ( .A(\align/N48 ), .B(sel_P[44]), .S0(n516), .Y(ali_P[44]) );
  MX2X1 U1349 ( .A(\align/N35 ), .B(sel_P[31]), .S0(n1030), .Y(ali_P[31]) );
  MX2X1 U1350 ( .A(\align/N33 ), .B(sel_P[29]), .S0(n1030), .Y(ali_P[29]) );
  MX2X1 U1351 ( .A(\align/N31 ), .B(sel_P[27]), .S0(n516), .Y(ali_P[27]) );
  MX2X1 U1352 ( .A(\align/N49 ), .B(sel_P[45]), .S0(n516), .Y(ali_P[45]) );
  MX2X1 U1353 ( .A(\align/N34 ), .B(sel_P[30]), .S0(n1030), .Y(ali_P[30]) );
  MX2X1 U1354 ( .A(\align/N51 ), .B(sel_P[47]), .S0(n516), .Y(ali_P[47]) );
  MX2X1 U1355 ( .A(\align/N50 ), .B(sel_P[46]), .S0(n516), .Y(ali_P[46]) );
  MX2X1 U1356 ( .A(\align/N32 ), .B(sel_P[28]), .S0(n516), .Y(ali_P[28]) );
  MXI2X1 U1357 ( .A(\align/sra_10/n188 ), .B(\align/sra_10/n192 ), .S0(n505), 
        .Y(\align/sra_10/n138 ) );
  MXI2X1 U1358 ( .A(\align/sra_10/n190 ), .B(\align/sra_10/n194 ), .S0(n505), 
        .Y(\align/sra_10/n140 ) );
  MXI2X1 U1359 ( .A(\align/sra_10/n199 ), .B(n508), .S0(n505), .Y(
        \align/sra_10/n149 ) );
  MXI2X1 U1360 ( .A(\align/sra_10/n200 ), .B(n508), .S0(n505), .Y(
        \align/sra_10/n150 ) );
  MXI2X1 U1361 ( .A(\align/sra_10/n198 ), .B(n508), .S0(n505), .Y(
        \align/sra_10/n148 ) );
  ADDFHX2 U1362 ( .A(\mul/mult_6/n191 ), .B(\mul/mult_6/n194 ), .CI(
        \mul/mult_6/n132 ), .CO(\mul/mult_6/n131 ), .S(sig_P[43]) );
  ADDFHX2 U1363 ( .A(\mul/mult_6/n216 ), .B(\mul/mult_6/n221 ), .CI(
        \mul/mult_6/n137 ), .CO(\mul/mult_6/n136 ), .S(sig_P[38]) );
  ADDFHX2 U1364 ( .A(\mul/mult_6/n222 ), .B(\mul/mult_6/n228 ), .CI(
        \mul/mult_6/n138 ), .CO(\mul/mult_6/n137 ), .S(sig_P[37]) );
  ADDFHX2 U1365 ( .A(\mul/mult_6/n236 ), .B(\mul/mult_6/n243 ), .CI(
        \mul/mult_6/n140 ), .CO(\mul/mult_6/n139 ), .S(sig_P[35]) );
  ADDFHX2 U1366 ( .A(\mul/mult_6/n244 ), .B(\mul/mult_6/n252 ), .CI(
        \mul/mult_6/n141 ), .CO(\mul/mult_6/n140 ), .S(sig_P[34]) );
  ADDFHX2 U1367 ( .A(\mul/mult_6/n262 ), .B(\mul/mult_6/n270 ), .CI(
        \mul/mult_6/n143 ), .CO(\mul/mult_6/n142 ), .S(sig_P[32]) );
  ADDFHX2 U1368 ( .A(\mul/mult_6/n379 ), .B(\mul/mult_6/n389 ), .CI(
        \mul/mult_6/n154 ), .CO(\mul/mult_6/n153 ), .S(sig_P[21]) );
  NAND2XL U1369 ( .A(\selc/N126 ), .B(n724), .Y(n762) );
  ADDFX2 U1370 ( .A(\mul/mult_6/n444 ), .B(\mul/mult_6/n450 ), .CI(
        \mul/mult_6/n161 ), .CO(\mul/mult_6/n160 ), .S(sig_P[14]) );
  ADDFX2 U1371 ( .A(\mul/mult_6/n451 ), .B(\mul/mult_6/n457 ), .CI(
        \mul/mult_6/n162 ), .CO(\mul/mult_6/n161 ), .S(sig_P[13]) );
  BUFX10 U1372 ( .A(n511), .Y(n505) );
  NAND2XL U1373 ( .A(\selc/N118 ), .B(n502), .Y(n770) );
  BUFX14 U1374 ( .A(sub_out[3]), .Y(n506) );
  BUFX8 U1375 ( .A(sub_out[3]), .Y(n705) );
  CMPR42X1 U1376 ( .A(\mul/mult_6/n297 ), .B(\mul/mult_6/n307 ), .C(
        \mul/mult_6/n294 ), .D(\mul/mult_6/n304 ), .ICI(\mul/mult_6/n300 ), 
        .S(\mul/mult_6/n291 ), .ICO(\mul/mult_6/n289 ), .CO(\mul/mult_6/n290 )
         );
  CMPR42X1 U1377 ( .A(\mul/mult_6/n817 ), .B(\mul/mult_6/n267 ), .C(
        \mul/mult_6/n256 ), .D(\mul/mult_6/n264 ), .ICI(\mul/mult_6/n260 ), 
        .S(\mul/mult_6/n253 ), .ICO(\mul/mult_6/n251 ), .CO(\mul/mult_6/n252 )
         );
  NAND2XL U1378 ( .A(\selc/N114 ), .B(n502), .Y(n774) );
  CMPR42X1 U1379 ( .A(\mul/mult_6/n405 ), .B(\mul/mult_6/n855 ), .C(
        \mul/mult_6/n831 ), .D(\mul/mult_6/n903 ), .ICI(\mul/mult_6/n411 ), 
        .S(\mul/mult_6/n403 ), .ICO(\mul/mult_6/n401 ), .CO(\mul/mult_6/n402 )
         );
  CMPR42X1 U1380 ( .A(\mul/mult_6/n876 ), .B(\mul/mult_6/n852 ), .C(
        \mul/mult_6/n384 ), .D(\mul/mult_6/n924 ), .ICI(\mul/mult_6/n380 ), 
        .S(\mul/mult_6/n371 ), .ICO(\mul/mult_6/n369 ), .CO(\mul/mult_6/n370 )
         );
  CMPR42X1 U1381 ( .A(\mul/mult_6/n376 ), .B(\mul/mult_6/n780 ), .C(
        \mul/mult_6/n383 ), .D(\mul/mult_6/n828 ), .ICI(\mul/mult_6/n804 ), 
        .S(\mul/mult_6/n374 ), .ICO(\mul/mult_6/n372 ), .CO(\mul/mult_6/n373 )
         );
  CMPR42X1 U1382 ( .A(\mul/mult_6/n387 ), .B(\mul/mult_6/n781 ), .C(
        \mul/mult_6/n396 ), .D(\mul/mult_6/n805 ), .ICI(\mul/mult_6/n829 ), 
        .S(\mul/mult_6/n385 ), .ICO(\mul/mult_6/n383 ), .CO(\mul/mult_6/n384 )
         );
  NAND2X2 U1383 ( .A(n689), .B(sig_B[0]), .Y(n536) );
  AOI22XL U1384 ( .A0(n700), .A1(sig_B[0]), .B0(n681), .B1(sig_B[1]), .Y(n564)
         );
  AOI22XL U1385 ( .A0(n699), .A1(sig_B[0]), .B0(n683), .B1(sig_B[1]), .Y(n529)
         );
  NAND2X2 U1386 ( .A(n685), .B(sig_B[0]), .Y(n531) );
  NAND2X2 U1387 ( .A(n687), .B(sig_B[0]), .Y(n530) );
  OR2X1 U1388 ( .A(\expadd/add_0_root_sub_0_root_sub_8/n2 ), .B(exp_C[0]), .Y(
        n660) );
  NAND3X2 U1389 ( .A(exp_A[0]), .B(exp_A[1]), .C(exp_A[2]), .Y(n1055) );
  AOI21X4 U1390 ( .A0(\ctrl/sub_0_root_add_0_root_sub_16/n24 ), .A1(n555), 
        .B0(\ctrl/sub_0_root_add_0_root_sub_16/n21 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n19 ) );
  INVX2 U1391 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n23 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n21 ) );
  XOR2X1 U1392 ( .A(n1033), .B(mux_out[7]), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/A[7] ) );
  MX2X1 U1393 ( .A(\ctrl/N27 ), .B(\ctrl/N11 ), .S0(n1043), .Y(D[23]) );
  NAND2X8 U1394 ( .A(n1042), .B(mux_out[1]), .Y(n1041) );
  NAND2X4 U1395 ( .A(\round/r298/n41 ), .B(\round/r298/n63 ), .Y(
        \round/r298/n40 ) );
  NAND3X2 U1396 ( .A(n522), .B(n993), .C(n992), .Y(n1002) );
  NAND3X2 U1397 ( .A(n998), .B(n997), .C(n996), .Y(n1001) );
  AND2X2 U1398 ( .A(\normal/N24 ), .B(n1043), .Y(n989) );
  AND2X2 U1399 ( .A(n999), .B(\normal/N70 ), .Y(n1000) );
  OAI21X1 U1400 ( .A0(\normal/srl_15/A[10] ), .A1(\normal/srl_15/A[8] ), .B0(
        n923), .Y(n935) );
  OR3X2 U1401 ( .A(n959), .B(n892), .C(n879), .Y(zero_cnt[4]) );
  INVX2 U1402 ( .A(n867), .Y(n868) );
  OAI21X1 U1403 ( .A0(n980), .A1(n979), .B0(n978), .Y(n981) );
  NAND2X2 U1404 ( .A(n875), .B(\normal/srl_15/A[21] ), .Y(n896) );
  AND2X8 U1405 ( .A(n887), .B(n889), .Y(n875) );
  AOI21X1 U1406 ( .A0(n977), .A1(n976), .B0(n975), .Y(n978) );
  INVX1 U1407 ( .A(n913), .Y(n930) );
  NOR2X2 U1408 ( .A(n877), .B(add_out[30]), .Y(n977) );
  OAI21XL U1409 ( .A0(\normal/srl_15/A[40] ), .A1(add_out[42]), .B0(n925), .Y(
        n926) );
  NAND2X2 U1410 ( .A(n869), .B(n842), .Y(n843) );
  NAND2X2 U1411 ( .A(n840), .B(n839), .Y(n874) );
  NAND2BX2 U1412 ( .AN(\normal/srl_15/A[32] ), .B(n837), .Y(n943) );
  INVXL U1413 ( .A(\normal/srl_15/A[21] ), .Y(n871) );
  OR2X2 U1414 ( .A(add_out[13]), .B(\normal/srl_15/A[11] ), .Y(n847) );
  OAI21X4 U1415 ( .A0(n501), .A1(n631), .B0(n815), .Y(add_out[19]) );
  AND2X4 U1416 ( .A(\sigadd/N51 ), .B(D[31]), .Y(add_out[49]) );
  INVXL U1417 ( .A(\normal/srl_15/A[44] ), .Y(n971) );
  INVX2 U1418 ( .A(add_out[31]), .Y(n837) );
  OAI21X4 U1419 ( .A0(n501), .A1(n620), .B0(n812), .Y(\normal/srl_15/A[22] )
         );
  OR2X2 U1420 ( .A(\normal/srl_15/A[44] ), .B(add_out[43]), .Y(n944) );
  OR2X2 U1421 ( .A(add_out[3]), .B(\normal/srl_15/A[4] ), .Y(n850) );
  OAI21X4 U1422 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n580), .B0(n792), .Y(
        add_out[42]) );
  XOR2X1 U1423 ( .A(\sigadd/sub_add_11_b0/n1 ), .B(n661), .Y(\sigadd/N51 ) );
  NAND2X2 U1424 ( .A(\sigadd/N43 ), .B(D[31]), .Y(n793) );
  NAND2X2 U1425 ( .A(\sigadd/N44 ), .B(D[31]), .Y(n792) );
  ADDHX1 U1426 ( .A(n620), .B(\sigadd/sub_add_11_b0/n28 ), .CO(
        \sigadd/sub_add_11_b0/n27 ), .S(\sigadd/N24 ) );
  ADDHX1 U1427 ( .A(n630), .B(\sigadd/sub_add_11_b0/n29 ), .CO(
        \sigadd/sub_add_11_b0/n28 ), .S(\sigadd/N23 ) );
  ADDHX1 U1428 ( .A(n621), .B(\sigadd/sub_add_11_b0/n30 ), .CO(
        \sigadd/sub_add_11_b0/n29 ), .S(\sigadd/N22 ) );
  ADDHX1 U1429 ( .A(n622), .B(\sigadd/sub_add_11_b0/n32 ), .CO(
        \sigadd/sub_add_11_b0/n31 ), .S(\sigadd/N20 ) );
  NAND2X2 U1430 ( .A(ali_P[0]), .B(ali_C[0]), .Y(\sigadd/add_9/n246 ) );
  OR2X2 U1431 ( .A(ali_P[32]), .B(ali_C[32]), .Y(n598) );
  OR2X2 U1432 ( .A(ali_P[34]), .B(ali_C[34]), .Y(n597) );
  OR2X2 U1433 ( .A(ali_P[36]), .B(ali_C[36]), .Y(n596) );
  OR2X2 U1434 ( .A(ali_P[38]), .B(ali_C[38]), .Y(n595) );
  MX2X1 U1435 ( .A(\align/N42 ), .B(sel_P[38]), .S0(n1030), .Y(ali_P[38]) );
  MX2X1 U1436 ( .A(\align/N46 ), .B(sel_P[42]), .S0(n1030), .Y(ali_P[42]) );
  MX2X1 U1437 ( .A(\align/N44 ), .B(sel_P[40]), .S0(n1030), .Y(ali_P[40]) );
  MX2X1 U1438 ( .A(\align/N41 ), .B(sel_P[37]), .S0(n1030), .Y(ali_P[37]) );
  MX2X1 U1439 ( .A(\align/N40 ), .B(sel_P[36]), .S0(n1030), .Y(ali_P[36]) );
  MX2X1 U1440 ( .A(\align/N45 ), .B(sel_P[41]), .S0(n1030), .Y(ali_P[41]) );
  MX2X1 U1441 ( .A(\align/N43 ), .B(sel_P[39]), .S0(n1030), .Y(ali_P[39]) );
  ADDFHX2 U1442 ( .A(\mul/mult_6/n335 ), .B(\mul/mult_6/n345 ), .CI(
        \mul/mult_6/n150 ), .CO(\mul/mult_6/n149 ), .S(sig_P[25]) );
  ADDFHX2 U1443 ( .A(\mul/mult_6/n357 ), .B(\mul/mult_6/n367 ), .CI(
        \mul/mult_6/n152 ), .CO(\mul/mult_6/n151 ), .S(sig_P[23]) );
  ADDFX2 U1444 ( .A(\mul/mult_6/n436 ), .B(\mul/mult_6/n443 ), .CI(
        \mul/mult_6/n160 ), .CO(\mul/mult_6/n159 ), .S(sig_P[15]) );
  NAND2XL U1445 ( .A(\selc/N117 ), .B(n502), .Y(n771) );
  BUFX20 U1446 ( .A(sub_out[0]), .Y(n507) );
  ADDFX1 U1447 ( .A(\mul/mult_6/n940 ), .B(\mul/mult_6/n487 ), .CI(
        \mul/mult_6/n169 ), .CO(\mul/mult_6/n168 ), .S(sig_P[6]) );
  INVX2 U1448 ( .A(n787), .Y(n517) );
  NAND2X2 U1449 ( .A(n787), .B(\two_en[1] ), .Y(n786) );
  ADDFX1 U1450 ( .A(\mul/mult_6/n941 ), .B(\mul/mult_6/n491 ), .CI(
        \mul/mult_6/n170 ), .CO(\mul/mult_6/n169 ), .S(sig_P[5]) );
  CMPR42X1 U1451 ( .A(\mul/mult_6/n764 ), .B(\mul/mult_6/n788 ), .C(
        \mul/mult_6/n224 ), .D(\mul/mult_6/n219 ), .ICI(\mul/mult_6/n220 ), 
        .S(\mul/mult_6/n216 ), .ICO(\mul/mult_6/n214 ), .CO(\mul/mult_6/n215 )
         );
  NAND2XL U1452 ( .A(\selc/N115 ), .B(n502), .Y(n773) );
  CMPR42X1 U1453 ( .A(\mul/mult_6/n201 ), .B(n650), .C(\mul/mult_6/n761 ), .D(
        \mul/mult_6/n205 ), .ICI(\mul/mult_6/n202 ), .S(\mul/mult_6/n199 ), 
        .ICO(\mul/mult_6/n197 ), .CO(\mul/mult_6/n198 ) );
  CMPR42X1 U1454 ( .A(\mul/mult_6/n275 ), .B(\mul/mult_6/n818 ), .C(
        \mul/mult_6/n794 ), .D(\mul/mult_6/n842 ), .ICI(\mul/mult_6/n268 ), 
        .S(\mul/mult_6/n265 ), .ICO(\mul/mult_6/n263 ), .CO(\mul/mult_6/n264 )
         );
  CMPR42X1 U1455 ( .A(\mul/mult_6/n820 ), .B(\mul/mult_6/n796 ), .C(
        \mul/mult_6/n295 ), .D(\mul/mult_6/n844 ), .ICI(\mul/mult_6/n296 ), 
        .S(\mul/mult_6/n284 ), .ICO(\mul/mult_6/n282 ), .CO(\mul/mult_6/n283 )
         );
  CMPR42X1 U1456 ( .A(\mul/mult_6/n867 ), .B(\mul/mult_6/n771 ), .C(
        \mul/mult_6/n819 ), .D(\mul/mult_6/n843 ), .ICI(\mul/mult_6/n277 ), 
        .S(\mul/mult_6/n274 ), .ICO(\mul/mult_6/n272 ), .CO(\mul/mult_6/n273 )
         );
  ADDFX1 U1457 ( .A(\mul/mult_6/n942 ), .B(\mul/mult_6/n493 ), .CI(
        \mul/mult_6/n171 ), .CO(\mul/mult_6/n170 ), .S(sig_P[4]) );
  CMPR42X1 U1458 ( .A(\mul/mult_6/n799 ), .B(\mul/mult_6/n328 ), .C(
        \mul/mult_6/n847 ), .D(\mul/mult_6/n871 ), .ICI(\mul/mult_6/n329 ), 
        .S(\mul/mult_6/n316 ), .ICO(\mul/mult_6/n314 ), .CO(\mul/mult_6/n315 )
         );
  CMPR42X1 U1459 ( .A(\mul/mult_6/n342 ), .B(\mul/mult_6/n776 ), .C(
        \mul/mult_6/n332 ), .D(\mul/mult_6/n824 ), .ICI(\mul/mult_6/n872 ), 
        .S(\mul/mult_6/n330 ), .ICO(\mul/mult_6/n328 ), .CO(\mul/mult_6/n329 )
         );
  CMPR42X1 U1460 ( .A(n674), .B(\mul/mult_6/n240 ), .C(n641), .D(
        \mul/mult_6/n814 ), .ICI(\mul/mult_6/n766 ), .S(\mul/mult_6/n232 ), 
        .ICO(\mul/mult_6/n230 ), .CO(\mul/mult_6/n231 ) );
  ADDFX1 U1461 ( .A(\mul/mult_6/n943 ), .B(\mul/mult_6/n495 ), .CI(
        \mul/mult_6/n172 ), .CO(\mul/mult_6/n171 ), .S(sig_P[3]) );
  CMPR42X1 U1462 ( .A(\mul/mult_6/n257 ), .B(n638), .C(\mul/mult_6/n840 ), .D(
        \mul/mult_6/n249 ), .ICI(\mul/mult_6/n254 ), .S(\mul/mult_6/n247 ), 
        .ICO(\mul/mult_6/n245 ), .CO(\mul/mult_6/n246 ) );
  ADDFX1 U1463 ( .A(\mul/mult_6/n489 ), .B(\mul/mult_6/n916 ), .CI(
        \mul/mult_6/n490 ), .CO(\mul/mult_6/n486 ), .S(\mul/mult_6/n487 ) );
  INVX2 U1464 ( .A(\mul/mult_6/n175 ), .Y(\mul/mult_6/n176 ) );
  ADDFX1 U1465 ( .A(\expadd/N4 ), .B(exp_B[4]), .CI(
        \expadd/add_0_root_sub_0_root_sub_8/n6 ), .CO(
        \expadd/add_0_root_sub_0_root_sub_8/n5 ), .S(exp_P[4]) );
  OA21X1 U1466 ( .A0(n1059), .A1(exp_A[6]), .B0(n1060), .Y(\expadd/N6 ) );
  NAND2BX8 U1467 ( .AN(\mul/mult_6/n1439 ), .B(\mul/mult_6/n1455 ), .Y(
        \mul/mult_6/n48 ) );
  NAND2BX8 U1468 ( .AN(\mul/mult_6/n1443 ), .B(\mul/mult_6/n1459 ), .Y(
        \mul/mult_6/n8 ) );
  NAND2X2 U1469 ( .A(n1056), .B(exp_A[4]), .Y(n1058) );
  OR2X2 U1470 ( .A(sig_B[21]), .B(sig_B[22]), .Y(n592) );
  INVX2 U1471 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n8 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n36 ) );
  OR2X2 U1472 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/A[4] ), .B(n708), .Y(
        n555) );
  INVX2 U1473 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n31 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n29 ) );
  OR2X2 U1474 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/A[2] ), .B(n712), .Y(
        n554) );
  OA21X4 U1475 ( .A0(n1042), .A1(mux_out[1]), .B0(n1041), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/A[1] ) );
  INVX2 U1476 ( .A(n1018), .Y(D[11]) );
  INVX2 U1477 ( .A(n1017), .Y(D[10]) );
  INVX2 U1478 ( .A(n1009), .Y(D[2]) );
  INVX2 U1479 ( .A(n1020), .Y(D[13]) );
  INVX2 U1480 ( .A(n1014), .Y(D[7]) );
  INVX2 U1481 ( .A(n1023), .Y(D[16]) );
  INVX2 U1482 ( .A(n1008), .Y(D[1]) );
  INVX2 U1483 ( .A(n1013), .Y(D[6]) );
  INVX2 U1484 ( .A(n1024), .Y(D[17]) );
  INVX2 U1485 ( .A(n1010), .Y(D[3]) );
  INVX2 U1486 ( .A(n1022), .Y(D[15]) );
  INVX2 U1487 ( .A(n1021), .Y(D[14]) );
  CLKXOR2X4 U1488 ( .A(n39), .B(\ctrl/add_1_root_add_16_2/A[0] ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/A[0] ) );
  INVXL U1489 ( .A(\round/r298/n52 ), .Y(\round/r298/n53 ) );
  NAND2X2 U1490 ( .A(\normal/N71 ), .B(n999), .Y(n987) );
  INVX2 U1491 ( .A(n503), .Y(n711) );
  OR2X6 U1492 ( .A(n966), .B(n965), .Y(zero_cnt[1]) );
  OR2X2 U1493 ( .A(n703), .B(\ctrl/add_1_root_add_16_2/A[4] ), .Y(n533) );
  AOI211X2 U1494 ( .A0(n916), .A1(add_out[17]), .B0(n915), .C0(n914), .Y(n917)
         );
  NAND2X2 U1495 ( .A(n868), .B(add_out[15]), .Y(n885) );
  NAND2XL U1496 ( .A(n875), .B(add_out[18]), .Y(n872) );
  NAND2X2 U1497 ( .A(n977), .B(n969), .Y(n956) );
  INVXL U1498 ( .A(n909), .Y(n910) );
  INVXL U1499 ( .A(n924), .Y(n925) );
  NAND2X8 U1500 ( .A(n832), .B(n972), .Y(n1043) );
  NAND2BX2 U1501 ( .AN(\normal/srl_15/A[8] ), .B(n849), .Y(n858) );
  INVXL U1502 ( .A(add_out[24]), .Y(n907) );
  NOR2X2 U1503 ( .A(\normal/srl_15/A[29] ), .B(add_out[26]), .Y(n840) );
  NOR2X2 U1504 ( .A(\normal/srl_15/A[9] ), .B(\normal/srl_15/A[6] ), .Y(n849)
         );
  OAI21X4 U1505 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n636), .B0(n826), .Y(
        \normal/srl_15/A[8] ) );
  OAI21X4 U1506 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n635), .B0(n824), .Y(
        \normal/srl_15/A[10] ) );
  INVXL U1507 ( .A(add_out[45]), .Y(n945) );
  NOR2X2 U1508 ( .A(add_out[30]), .B(add_out[28]), .Y(n839) );
  INVXL U1509 ( .A(\normal/srl_15/A[40] ), .Y(n908) );
  INVX2 U1510 ( .A(\normal/srl_15/A[32] ), .Y(n884) );
  OAI21X1 U1511 ( .A0(n895), .A1(\normal/srl_15/A[4] ), .B0(n894), .Y(n900) );
  INVXL U1512 ( .A(\normal/srl_15/A[1] ), .Y(n851) );
  NAND2X2 U1513 ( .A(\sigadd/N16 ), .B(n501), .Y(n820) );
  NAND2X2 U1514 ( .A(\sigadd/N20 ), .B(n501), .Y(n816) );
  NAND2X2 U1515 ( .A(\sigadd/N24 ), .B(n501), .Y(n812) );
  ADDHX1 U1516 ( .A(n632), .B(\sigadd/sub_add_11_b0/n33 ), .CO(
        \sigadd/sub_add_11_b0/n32 ), .S(\sigadd/N19 ) );
  ADDHX1 U1517 ( .A(n646), .B(\sigadd/sub_add_11_b0/n39 ), .CO(
        \sigadd/sub_add_11_b0/n38 ), .S(\sigadd/N13 ) );
  INVXL U1518 ( .A(\sigadd/add_9/n235 ), .Y(\sigadd/add_9/n293 ) );
  INVXL U1519 ( .A(\sigadd/add_9/n243 ), .Y(\sigadd/add_9/n295 ) );
  INVX2 U1520 ( .A(\sigadd/add_9/n209 ), .Y(\sigadd/add_9/n207 ) );
  INVXL U1521 ( .A(\sigadd/add_9/n227 ), .Y(\sigadd/add_9/n291 ) );
  INVXL U1522 ( .A(\sigadd/add_9/n219 ), .Y(\sigadd/add_9/n289 ) );
  INVXL U1523 ( .A(\sigadd/add_9/n211 ), .Y(\sigadd/add_9/n287 ) );
  OR2X2 U1524 ( .A(ali_P[28]), .B(ali_C[28]), .Y(n573) );
  OR2X2 U1525 ( .A(ali_P[18]), .B(ali_C[18]), .Y(n578) );
  OR2X2 U1526 ( .A(ali_P[16]), .B(ali_C[16]), .Y(n579) );
  OR2X2 U1527 ( .A(ali_P[22]), .B(ali_C[22]), .Y(n576) );
  OR2X2 U1528 ( .A(ali_P[24]), .B(ali_C[24]), .Y(n575) );
  OR2X2 U1529 ( .A(ali_P[20]), .B(ali_C[20]), .Y(n577) );
  OR2X2 U1530 ( .A(ali_P[26]), .B(ali_C[26]), .Y(n574) );
  OR2X2 U1531 ( .A(ali_P[30]), .B(ali_C[30]), .Y(n599) );
  INVX2 U1532 ( .A(sig_P[41]), .Y(\selc/r299/A[41] ) );
  NAND2XL U1533 ( .A(n719), .B(n716), .Y(\align/sra_11/n754 ) );
  NAND2XL U1534 ( .A(\selc/N124 ), .B(n724), .Y(n764) );
  NAND2XL U1535 ( .A(\selc/N123 ), .B(n724), .Y(n765) );
  NAND2XL U1536 ( .A(n506), .B(\align/sra_11/n624 ), .Y(\align/sra_11/n697 )
         );
  NAND2XL U1537 ( .A(n506), .B(\align/sra_11/n630 ), .Y(\align/sra_11/n718 )
         );
  NAND2XL U1538 ( .A(\selc/N122 ), .B(n724), .Y(n766) );
  NAND2XL U1539 ( .A(n506), .B(\align/sra_11/n618 ), .Y(\align/sra_11/n684 )
         );
  NAND2XL U1540 ( .A(n506), .B(\align/sra_11/n612 ), .Y(\align/sra_11/n672 )
         );
  NAND2XL U1541 ( .A(n506), .B(\align/sra_11/n471 ), .Y(\align/sra_11/n468 )
         );
  NAND2XL U1542 ( .A(n506), .B(\align/sra_11/n652 ), .Y(\align/sra_11/n736 )
         );
  NAND2XL U1543 ( .A(n506), .B(\align/sra_11/n646 ), .Y(\align/sra_11/n729 )
         );
  NAND2XL U1544 ( .A(n506), .B(\align/sra_11/n478 ), .Y(\align/sra_11/n475 )
         );
  NAND2XL U1545 ( .A(\selc/N121 ), .B(n724), .Y(n767) );
  NAND2X1 U1546 ( .A(\align/sra_11/SH[1] ), .B(n653), .Y(\align/sra_11/n723 )
         );
  NAND2X1 U1547 ( .A(\align/sra_11/SH[1] ), .B(\align/sra_11/n709 ), .Y(
        \align/sra_11/n663 ) );
  NAND2XL U1548 ( .A(\selc/N120 ), .B(n724), .Y(n768) );
  AND2X1 U1549 ( .A(n507), .B(sel_C[23]), .Y(n653) );
  NAND2XL U1550 ( .A(\selc/N119 ), .B(n724), .Y(n769) );
  BUFX10 U1551 ( .A(sub_out[4]), .Y(n719) );
  BUFX12 U1552 ( .A(\align/sra_11/n465 ), .Y(n510) );
  MX2X4 U1553 ( .A(\sub/N17 ), .B(\sub/N8 ), .S0(n516), .Y(sub_out[3]) );
  NAND2XL U1554 ( .A(\selc/N116 ), .B(n502), .Y(n772) );
  INVX2 U1555 ( .A(n780), .Y(n785) );
  OAI21X1 U1556 ( .A0(exp_C[6]), .A1(n1031), .B0(n779), .Y(n781) );
  NAND2BX2 U1557 ( .AN(exp_P[7]), .B(exp_C[7]), .Y(n780) );
  INVX2 U1558 ( .A(exp_P[6]), .Y(n1031) );
  OA22X2 U1559 ( .A0(exp_P[6]), .A1(n1032), .B0(exp_P[5]), .B1(n1029), .Y(n778) );
  INVX2 U1560 ( .A(\mul/mult_6/n580 ), .Y(\mul/mult_6/n575 ) );
  XOR2X1 U1561 ( .A(exp_A[7]), .B(n1060), .Y(
        \expadd/add_0_root_sub_0_root_sub_8/B[7] ) );
  CLKNAND2X2 U1562 ( .A(n679), .B(sig_B[0]), .Y(n524) );
  NAND2X2 U1563 ( .A(n692), .B(sig_B[0]), .Y(n586) );
  AOI21X1 U1564 ( .A0(n1058), .A1(n1057), .B0(n1059), .Y(\expadd/N5 ) );
  NAND2X2 U1565 ( .A(n1059), .B(exp_A[6]), .Y(n1060) );
  INVX2 U1566 ( .A(\mul/mult_6/n608 ), .Y(\mul/mult_6/n715 ) );
  NAND2BX8 U1567 ( .AN(\mul/mult_6/n1441 ), .B(\mul/mult_6/n1457 ), .Y(
        \mul/mult_6/n28 ) );
  NAND2BX8 U1568 ( .AN(\mul/mult_6/n1442 ), .B(\mul/mult_6/n1458 ), .Y(
        \mul/mult_6/n18 ) );
  NOR2X4 U1569 ( .A(\mul/mult_6/n1442 ), .B(\mul/mult_6/n1458 ), .Y(
        \mul/mult_6/n12 ) );
  NOR2X4 U1570 ( .A(\mul/mult_6/n1459 ), .B(\mul/mult_6/n1443 ), .Y(
        \mul/mult_6/n2 ) );
  INVX2 U1571 ( .A(\mul/mult_6/n705 ), .Y(\mul/mult_6/n731 ) );
  INVX2 U1572 ( .A(\mul/mult_6/n697 ), .Y(\mul/mult_6/n695 ) );
  INVX2 U1573 ( .A(\mul/mult_6/n691 ), .Y(\mul/mult_6/n728 ) );
  INVX2 U1574 ( .A(\mul/mult_6/n686 ), .Y(\mul/mult_6/n727 ) );
  INVX2 U1575 ( .A(exp_A[3]), .Y(n1054) );
  INVX2 U1576 ( .A(exp_A[5]), .Y(n1057) );
  AOI21X4 U1577 ( .A0(\ctrl/sub_0_root_add_0_root_sub_16/n32 ), .A1(n554), 
        .B0(\ctrl/sub_0_root_add_0_root_sub_16/n29 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n27 ) );
  AND2X2 U1578 ( .A(\ctrl/add_1_root_add_16_2/n17 ), .B(
        \ctrl/add_1_root_add_16_2/n13 ), .Y(n585) );
  AND2X2 U1579 ( .A(\ctrl/add_1_root_add_16_2/n16 ), .B(
        \ctrl/add_1_root_add_16_2/n13 ), .Y(n526) );
  NOR2X2 U1580 ( .A(n995), .B(n994), .Y(n996) );
  INVX2 U1581 ( .A(\ctrl/add_1_root_add_16_2/n62 ), .Y(
        \ctrl/add_1_root_add_16_2/n60 ) );
  NAND2X2 U1582 ( .A(n503), .B(\ctrl/add_1_root_add_16_2/A[0] ), .Y(
        \ctrl/add_1_root_add_16_2/n62 ) );
  INVX2 U1583 ( .A(n504), .Y(n713) );
  INVX2 U1584 ( .A(n512), .Y(n712) );
  INVX2 U1585 ( .A(n513), .Y(n709) );
  NAND2X2 U1586 ( .A(n715), .B(mux_out[1]), .Y(\ctrl/add_1_root_add_16_2/n57 )
         );
  INVX2 U1587 ( .A(n715), .Y(n710) );
  INVX2 U1588 ( .A(n703), .Y(n708) );
  NAND2BX8 U1589 ( .AN(n897), .B(n835), .Y(n941) );
  INVXL U1590 ( .A(n858), .Y(n862) );
  INVXL U1591 ( .A(n874), .Y(n878) );
  OAI21X4 U1592 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n647), .B0(n825), .Y(
        \normal/srl_15/A[9] ) );
  AOI2B1X1 U1593 ( .A1N(\normal/srl_15/A[36] ), .A0(add_out[35]), .B0(
        add_out[37]), .Y(n898) );
  OAI21X4 U1594 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n623), .B0(n818), .Y(
        add_out[16]) );
  OAI21X4 U1595 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n632), .B0(n817), .Y(
        add_out[17]) );
  OAI21X4 U1596 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n614), .B0(n807), .Y(
        \normal/srl_15/A[27] ) );
  INVX2 U1597 ( .A(add_out[2]), .Y(n866) );
  ADDHX2 U1598 ( .A(n560), .B(\sigadd/sub_add_11_b0/n2 ), .CO(
        \sigadd/sub_add_11_b0/n1 ), .S(\sigadd/N50 ) );
  ADDHX2 U1599 ( .A(n568), .B(\sigadd/sub_add_11_b0/n3 ), .CO(
        \sigadd/sub_add_11_b0/n2 ), .S(\sigadd/N49 ) );
  ADDHX2 U1600 ( .A(n558), .B(\sigadd/sub_add_11_b0/n4 ), .CO(
        \sigadd/sub_add_11_b0/n3 ), .S(\sigadd/N48 ) );
  ADDHX2 U1601 ( .A(n588), .B(\sigadd/sub_add_11_b0/n11 ), .CO(
        \sigadd/sub_add_11_b0/n10 ), .S(\sigadd/N41 ) );
  ADDHX2 U1602 ( .A(n582), .B(\sigadd/sub_add_11_b0/n12 ), .CO(
        \sigadd/sub_add_11_b0/n11 ), .S(\sigadd/N40 ) );
  ADDHX2 U1603 ( .A(n611), .B(\sigadd/sub_add_11_b0/n17 ), .CO(
        \sigadd/sub_add_11_b0/n16 ), .S(\sigadd/N35 ) );
  ADDHX2 U1604 ( .A(n600), .B(\sigadd/sub_add_11_b0/n18 ), .CO(
        \sigadd/sub_add_11_b0/n17 ), .S(\sigadd/N34 ) );
  ADDHX1 U1605 ( .A(n634), .B(\sigadd/sub_add_11_b0/n38 ), .CO(
        \sigadd/sub_add_11_b0/n37 ), .S(\sigadd/N14 ) );
  INVXL U1606 ( .A(\sigadd/add_9/n75 ), .Y(\sigadd/add_9/n253 ) );
  INVXL U1607 ( .A(\sigadd/add_9/n83 ), .Y(\sigadd/add_9/n255 ) );
  INVXL U1608 ( .A(\sigadd/add_9/n59 ), .Y(\sigadd/add_9/n249 ) );
  INVXL U1609 ( .A(\sigadd/add_9/n179 ), .Y(\sigadd/add_9/n279 ) );
  INVXL U1610 ( .A(\sigadd/add_9/n203 ), .Y(\sigadd/add_9/n285 ) );
  INVXL U1611 ( .A(\sigadd/add_9/n67 ), .Y(\sigadd/add_9/n251 ) );
  INVXL U1612 ( .A(\sigadd/add_9/n195 ), .Y(\sigadd/add_9/n283 ) );
  INVXL U1613 ( .A(\sigadd/add_9/n187 ), .Y(\sigadd/add_9/n281 ) );
  MXI2X2 U1614 ( .A(n1028), .B(n1045), .S0(n516), .Y(mux_out[1]) );
  BUFX20 U1615 ( .A(sub_out[1]), .Y(\align/sra_11/SH[1] ) );
  INVXL U1616 ( .A(exp_P[7]), .Y(\sub/sub_17/n10 ) );
  AOI22X2 U1617 ( .A0(n701), .A1(sig_B[0]), .B0(n679), .B1(sig_B[1]), .Y(n523)
         );
  INVX2 U1618 ( .A(\mul/mult_6/n653 ), .Y(\mul/mult_6/n655 ) );
  INVX2 U1619 ( .A(\mul/mult_6/n20 ), .Y(n682) );
  INVX2 U1620 ( .A(\mul/mult_6/n30 ), .Y(n684) );
  INVX2 U1621 ( .A(\mul/mult_6/n9 ), .Y(n680) );
  INVX2 U1622 ( .A(\mul/mult_6/n630 ), .Y(\mul/mult_6/n718 ) );
  NAND2BX8 U1623 ( .AN(\mul/mult_6/n1438 ), .B(\mul/mult_6/n1454 ), .Y(
        \mul/mult_6/n58 ) );
  NAND2BX8 U1624 ( .AN(\mul/mult_6/n1440 ), .B(\mul/mult_6/n1456 ), .Y(
        \mul/mult_6/n38 ) );
  NAND2BX8 U1625 ( .AN(\mul/mult_6/n1436 ), .B(\mul/mult_6/n1452 ), .Y(
        \mul/mult_6/n76 ) );
  NAND2BX8 U1626 ( .AN(\mul/mult_6/n1437 ), .B(\mul/mult_6/n1453 ), .Y(
        \mul/mult_6/n68 ) );
  NOR2X4 U1627 ( .A(\mul/mult_6/n1437 ), .B(\mul/mult_6/n1453 ), .Y(
        \mul/mult_6/n62 ) );
  INVX4 U1628 ( .A(\two_en[1] ), .Y(n722) );
  INVX4 U1629 ( .A(\two_en[1] ), .Y(n721) );
  OR2X2 U1630 ( .A(n503), .B(\ctrl/add_1_root_add_16_2/A[0] ), .Y(n520) );
  OR2X2 U1631 ( .A(n715), .B(mux_out[1]), .Y(n534) );
  MXI2X1 U1632 ( .A(\align/sra_10/n117 ), .B(\align/sra_10/n125 ), .S0(n506), 
        .Y(\align/sra_10/n67 ) );
  BUFX10 U1633 ( .A(n515), .Y(n717) );
  CLKAND2X12 U1634 ( .A(n783), .B(n782), .Y(n787) );
  ADDHX1 U1635 ( .A(n631), .B(\sigadd/sub_add_11_b0/n31 ), .CO(
        \sigadd/sub_add_11_b0/n30 ), .S(\sigadd/N21 ) );
  OAI21X4 U1636 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n645), .B0(n821), .Y(
        add_out[13]) );
  ADDHX1 U1637 ( .A(n645), .B(\sigadd/sub_add_11_b0/n37 ), .CO(
        \sigadd/sub_add_11_b0/n36 ), .S(\sigadd/N15 ) );
  INVX4 U1638 ( .A(\two_en[1] ), .Y(n723) );
  OAI21X8 U1639 ( .A0(n785), .A1(n784), .B0(n787), .Y(n1030) );
  NAND2BX8 U1640 ( .AN(n949), .B(n948), .Y(n897) );
  NOR2X8 U1641 ( .A(n924), .B(add_out[42]), .Y(n909) );
  NAND2BX8 U1642 ( .AN(n1043), .B(n833), .Y(n924) );
  OA21X1 U1643 ( .A0(\mul/mult_6/n1387 ), .A1(\mul/mult_6/n76 ), .B0(n538), 
        .Y(n609) );
  MXI2X2 U1644 ( .A(n1029), .B(n1047), .S0(n516), .Y(mux_out[5]) );
  NOR2X8 U1645 ( .A(n913), .B(n843), .Y(n887) );
  NAND2BX8 U1646 ( .AN(n942), .B(n838), .Y(n877) );
  INVXL U1647 ( .A(\sigadd/add_9/n171 ), .Y(\sigadd/add_9/n277 ) );
  INVXL U1648 ( .A(\sigadd/add_9/n163 ), .Y(\sigadd/add_9/n275 ) );
  INVXL U1649 ( .A(\sigadd/add_9/n155 ), .Y(\sigadd/add_9/n273 ) );
  INVXL U1650 ( .A(\sigadd/add_9/n147 ), .Y(\sigadd/add_9/n271 ) );
  CLKXOR2X2 U1651 ( .A(\mul/mult_6/n698 ), .B(\mul/mult_6/n570 ), .Y(n545) );
  OA21X1 U1652 ( .A0(\mul/mult_6/n1386 ), .A1(\mul/mult_6/n76 ), .B0(
        \mul/mult_6/n996 ), .Y(n608) );
  INVX2 U1653 ( .A(\mul/mult_6/n666 ), .Y(\mul/mult_6/n664 ) );
  INVXL U1654 ( .A(n941), .Y(n953) );
  INVXL U1655 ( .A(n859), .Y(n860) );
  NAND2X8 U1656 ( .A(n859), .B(n846), .Y(n968) );
  NAND2BX8 U1657 ( .AN(n980), .B(n979), .Y(n931) );
  NAND2BX8 U1658 ( .AN(n877), .B(n841), .Y(n913) );
  INVXL U1659 ( .A(\sigadd/add_9/n139 ), .Y(\sigadd/add_9/n269 ) );
  INVXL U1660 ( .A(\sigadd/add_9/n131 ), .Y(\sigadd/add_9/n267 ) );
  INVXL U1661 ( .A(\sigadd/add_9/n123 ), .Y(\sigadd/add_9/n265 ) );
  INVX2 U1662 ( .A(\mul/mult_6/n50 ), .Y(n688) );
  INVX2 U1663 ( .A(\mul/mult_6/n40 ), .Y(n686) );
  OA21X1 U1664 ( .A0(n546), .A1(\mul/mult_6/n76 ), .B0(\mul/mult_6/n995 ), .Y(
        n606) );
  INVX2 U1665 ( .A(\mul/mult_6/n652 ), .Y(\mul/mult_6/n654 ) );
  INVX2 U1666 ( .A(\mul/mult_6/n670 ), .Y(\mul/mult_6/n668 ) );
  MXI2X2 U1667 ( .A(n1049), .B(\sub/sub_17/n14 ), .S0(n516), .Y(mux_out[3]) );
  NOR2X8 U1668 ( .A(n867), .B(add_out[15]), .Y(n859) );
  NAND2BX8 U1669 ( .AN(n940), .B(n873), .Y(n867) );
  NAND2BX8 U1670 ( .AN(n941), .B(n836), .Y(n942) );
  INVXL U1671 ( .A(\sigadd/add_9/n115 ), .Y(\sigadd/add_9/n263 ) );
  INVXL U1672 ( .A(\sigadd/add_9/n107 ), .Y(\sigadd/add_9/n261 ) );
  OR2X2 U1673 ( .A(ali_P[48]), .B(ali_C[48]), .Y(n617) );
  INVX2 U1674 ( .A(\mul/mult_6/n665 ), .Y(\mul/mult_6/n723 ) );
  INVX2 U1675 ( .A(\mul/mult_6/n671 ), .Y(\mul/mult_6/n669 ) );
  INVXL U1676 ( .A(n887), .Y(n890) );
  NAND2BX8 U1677 ( .AN(n968), .B(n938), .Y(n853) );
  NAND2BX8 U1678 ( .AN(n931), .B(n845), .Y(n940) );
  OAI21X4 U1679 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n568), .B0(n830), .Y(
        add_out[47]) );
  OAI21X4 U1680 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n558), .B0(n788), .Y(
        add_out[46]) );
  INVXL U1681 ( .A(\sigadd/add_9/n99 ), .Y(\sigadd/add_9/n259 ) );
  INVXL U1682 ( .A(\sigadd/add_9/n91 ), .Y(\sigadd/add_9/n257 ) );
  OR2X2 U1683 ( .A(ali_P[46]), .B(ali_C[46]), .Y(n618) );
  NOR2BX1 U1684 ( .AN(exp_A[1]), .B(\expadd/add_0_root_sub_0_root_sub_8/B[0] ), 
        .Y(n1053) );
  INVX2 U1685 ( .A(exp_A[0]), .Y(\expadd/add_0_root_sub_0_root_sub_8/B[0] ) );
  INVX2 U1686 ( .A(\mul/mult_6/n620 ), .Y(\mul/mult_6/n717 ) );
  AOI21X4 U1687 ( .A0(n1034), .A1(n1035), .B0(n1033), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n10 ) );
  AOI21X4 U1688 ( .A0(n1037), .A1(n1038), .B0(n1036), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/A[4] ) );
  NOR2BX8 U1689 ( .AN(\ctrl/add_1_root_add_16_2/A[4] ), .B(n1038), .Y(n1036)
         );
  NAND2X8 U1690 ( .A(n901), .B(n894), .Y(n903) );
  NOR2X8 U1691 ( .A(n853), .B(n847), .Y(n923) );
  OAI21X4 U1692 ( .A0(n501), .A1(n616), .B0(n811), .Y(add_out[23]) );
  MX2X1 U1693 ( .A(\sub/N18 ), .B(\sub/N9 ), .S0(n516), .Y(sub_out[4]) );
  CLKINVX40 U1694 ( .A(n519), .Y(n707) );
  INVX2 U1695 ( .A(\mul/mult_6/n696 ), .Y(\mul/mult_6/n729 ) );
  INVX2 U1696 ( .A(\mul/mult_6/n387 ), .Y(\mul/mult_6/n386 ) );
  INVX2 U1697 ( .A(\mul/mult_6/n614 ), .Y(\mul/mult_6/n612 ) );
  INVX2 U1698 ( .A(\mul/mult_6/n613 ), .Y(\mul/mult_6/n611 ) );
  INVX2 U1699 ( .A(\mul/mult_6/n635 ), .Y(\mul/mult_6/n719 ) );
  INVX2 U1700 ( .A(\mul/mult_6/n649 ), .Y(\mul/mult_6/n721 ) );
  NOR2BX4 U1701 ( .AN(\ctrl/add_1_root_add_16_2/n13 ), .B(n1035), .Y(n1033) );
  OA21X4 U1702 ( .A0(n1039), .A1(mux_out[3]), .B0(n1038), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/A[3] ) );
  NAND2X8 U1703 ( .A(n923), .B(n848), .Y(n964) );
  OAI21X4 U1704 ( .A0(n501), .A1(n603), .B0(n808), .Y(add_out[26]) );
  OAI2BB1X1 U1705 ( .A0N(n517), .A1N(\align/N102 ), .B0(n786), .Y(ali_C[48])
         );
  OAI2BB1X1 U1706 ( .A0N(n517), .A1N(\align/N101 ), .B0(n786), .Y(ali_C[47])
         );
  OA21X1 U1707 ( .A0(n1053), .A1(exp_A[2]), .B0(n1055), .Y(\expadd/N2 ) );
  OA21X1 U1708 ( .A0(n1056), .A1(exp_A[4]), .B0(n1058), .Y(\expadd/N4 ) );
  INVX2 U1709 ( .A(\mul/mult_6/n596 ), .Y(\mul/mult_6/n713 ) );
  NAND2X2 U1710 ( .A(n695), .B(sig_B[0]), .Y(n537) );
  OA21X4 U1711 ( .A0(n1036), .A1(mux_out[5]), .B0(n1035), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/A[5] ) );
  NOR2X8 U1712 ( .A(n1041), .B(n1040), .Y(n1039) );
  AND2X8 U1713 ( .A(\round/r298/n1 ), .B(n563), .Y(n521) );
  NOR3X8 U1714 ( .A(n964), .B(add_out[7]), .C(n858), .Y(n901) );
  MX2X1 U1715 ( .A(\sub/N16 ), .B(\sub/N7 ), .S0(n516), .Y(sub_out[2]) );
  NAND3X2 U1716 ( .A(n920), .B(n918), .C(add_out[7]), .Y(n856) );
  OR2XL U1717 ( .A(\mul/mult_6/n946 ), .B(sig_A[2]), .Y(n640) );
  CLKAND2X12 U1718 ( .A(n521), .B(n1007), .Y(n39) );
  OAI21X4 U1719 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n581), .B0(n794), .Y(
        \normal/srl_15/A[40] ) );
  OAI21X4 U1720 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n566), .B0(n789), .Y(
        add_out[45]) );
  NOR2BX1 U1721 ( .AN(\align/N54 ), .B(n787), .Y(ali_C[0]) );
  INVX2 U1722 ( .A(exp_C[7]), .Y(n1027) );
  INVX2 U1723 ( .A(sig_A[17]), .Y(n664) );
  INVX2 U1724 ( .A(sig_B[13]), .Y(n673) );
  INVX2 U1725 ( .A(sig_B[12]), .Y(n674) );
  INVX2 U1726 ( .A(\mul/mult_6/n70 ), .Y(n694) );
  INVX2 U1727 ( .A(\mul/mult_6/n60 ), .Y(n691) );
  INVX2 U1728 ( .A(sig_B[6]), .Y(n677) );
  INVX2 U1729 ( .A(\mul/mult_6/n591 ), .Y(\mul/mult_6/n712 ) );
  INVX2 U1730 ( .A(\mul/mult_6/n597 ), .Y(\mul/mult_6/n595 ) );
  INVX2 U1731 ( .A(\mul/mult_6/n603 ), .Y(\mul/mult_6/n714 ) );
  INVX2 U1732 ( .A(\mul/mult_6/n609 ), .Y(\mul/mult_6/n607 ) );
  INVX2 U1733 ( .A(\mul/mult_6/n615 ), .Y(\mul/mult_6/n716 ) );
  INVX2 U1734 ( .A(\mul/mult_6/n621 ), .Y(\mul/mult_6/n619 ) );
  INVX2 U1735 ( .A(\mul/mult_6/n636 ), .Y(\mul/mult_6/n634 ) );
  INVX2 U1736 ( .A(\mul/mult_6/n644 ), .Y(\mul/mult_6/n720 ) );
  INVX2 U1737 ( .A(\mul/mult_6/n650 ), .Y(\mul/mult_6/n648 ) );
  INVX2 U1738 ( .A(\mul/mult_6/n660 ), .Y(\mul/mult_6/n722 ) );
  INVX2 U1739 ( .A(\mul/mult_6/n672 ), .Y(\mul/mult_6/n724 ) );
  NAND2X2 U1740 ( .A(n1025), .B(n522), .Y(n1006) );
  INVX2 U1741 ( .A(n1011), .Y(D[4]) );
  INVX2 U1742 ( .A(\round/r298/n113 ), .Y(\round/r298/n112 ) );
  INVX2 U1743 ( .A(n1015), .Y(D[8]) );
  INVX2 U1744 ( .A(n1016), .Y(D[9]) );
  INVX2 U1745 ( .A(n1019), .Y(D[12]) );
  INVX2 U1746 ( .A(norm_out[14]), .Y(\round/r298/n73 ) );
  INVX2 U1747 ( .A(norm_out[16]), .Y(\round/r298/n61 ) );
  INVX2 U1748 ( .A(\round/r298/n63 ), .Y(\round/r298/n64 ) );
  INVX2 U1749 ( .A(n1012), .Y(D[5]) );
  INVX2 U1750 ( .A(norm_out[8]), .Y(\round/r298/n103 ) );
  INVX2 U1751 ( .A(norm_out[22]), .Y(\round/r298/n28 ) );
  INVX2 U1752 ( .A(\round/r298/n18 ), .Y(\round/r298/n19 ) );
  INVX2 U1753 ( .A(norm_out[24]), .Y(\round/r298/n16 ) );
  INVX2 U1754 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n33 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n40 ) );
  INVX2 U1755 ( .A(\ctrl/add_1_root_add_16_2/n36 ), .Y(
        \ctrl/add_1_root_add_16_2/n67 ) );
  INVX2 U1756 ( .A(\ctrl/sub_0_root_add_0_root_sub_16/n25 ), .Y(
        \ctrl/sub_0_root_add_0_root_sub_16/n38 ) );
  NAND2BX2 U1757 ( .AN(exp_P[7]), .B(n1027), .Y(mux_out[7]) );
  INVX2 U1758 ( .A(\ctrl/add_1_root_add_16_2/n13 ), .Y(n1034) );
  INVX2 U1759 ( .A(\ctrl/add_1_root_add_16_2/n18 ), .Y(
        \ctrl/add_1_root_add_16_2/n65 ) );
  INVX2 U1760 ( .A(\ctrl/add_1_root_add_16_2/n24 ), .Y(
        \ctrl/add_1_root_add_16_2/n22 ) );
  INVX2 U1761 ( .A(\ctrl/add_1_root_add_16_2/n28 ), .Y(
        \ctrl/add_1_root_add_16_2/n26 ) );
  OR2X2 U1762 ( .A(\ctrl/add_1_root_add_16_2/n41 ), .B(
        \ctrl/add_1_root_add_16_2/n36 ), .Y(n525) );
  INVX2 U1763 ( .A(\ctrl/add_1_root_add_16_2/A[4] ), .Y(n1037) );
  OR2X2 U1764 ( .A(\normal/N66 ), .B(\normal/N67 ), .Y(n994) );
  OR3X2 U1765 ( .A(\normal/N68 ), .B(\normal/N69 ), .C(\normal/N49 ), .Y(n995)
         );
  NAND2X2 U1766 ( .A(\normal/N25 ), .B(n1043), .Y(n988) );
  AOI211X2 U1767 ( .A0(n930), .A1(add_out[24]), .B0(n929), .C0(n928), .Y(n934)
         );
  INVX2 U1768 ( .A(add_out[34]), .Y(n927) );
  INVX2 U1769 ( .A(add_out[3]), .Y(n895) );
  NOR4X2 U1770 ( .A(n893), .B(n915), .C(n892), .D(n891), .Y(n902) );
  NOR4X2 U1771 ( .A(n883), .B(n882), .C(\normal/srl_15/A[9] ), .D(add_out[7]), 
        .Y(n893) );
  INVX2 U1772 ( .A(\normal/srl_15/A[6] ), .Y(n882) );
  INVX2 U1773 ( .A(n920), .Y(n883) );
  INVX2 U1774 ( .A(\normal/srl_15/A[4] ), .Y(n904) );
  NOR2X2 U1775 ( .A(add_out[2]), .B(\sigadd/sig[0] ), .Y(n880) );
  NOR4X2 U1776 ( .A(n961), .B(n960), .C(n959), .D(n958), .Y(n962) );
  AOI211X2 U1777 ( .A0(n953), .A1(n952), .B0(n951), .C0(n950), .Y(n954) );
  OR2X2 U1778 ( .A(\normal/srl_15/A[36] ), .B(add_out[35]), .Y(n952) );
  INVX2 U1779 ( .A(add_out[28]), .Y(n957) );
  INVX2 U1780 ( .A(add_out[16]), .Y(n939) );
  INVX2 U1781 ( .A(\normal/srl_15/A[8] ), .Y(n963) );
  INVX2 U1782 ( .A(\normal/srl_15/A[29] ), .Y(n969) );
  INVX2 U1783 ( .A(\normal/srl_15/A[27] ), .Y(n970) );
  AOI211X2 U1784 ( .A0(n901), .A1(add_out[5]), .B0(n966), .C0(n863), .Y(n865)
         );
  NOR4X2 U1785 ( .A(add_out[14]), .B(\normal/srl_15/A[10] ), .C(
        \normal/srl_15/A[12] ), .D(add_out[13]), .Y(n861) );
  NAND2X2 U1786 ( .A(n982), .B(n854), .Y(n855) );
  INVX2 U1787 ( .A(add_out[13]), .Y(n854) );
  INVX2 U1788 ( .A(\normal/srl_15/A[11] ), .Y(n852) );
  INVX2 U1789 ( .A(\normal/srl_15/A[9] ), .Y(n918) );
  INVX2 U1790 ( .A(\sigadd/add_9/n50 ), .Y(\sigadd/sig[0] ) );
  INVX2 U1791 ( .A(\sigadd/N7 ), .Y(n829) );
  NAND2X2 U1792 ( .A(\sigadd/N21 ), .B(n501), .Y(n815) );
  NAND2X2 U1793 ( .A(\sigadd/N23 ), .B(n501), .Y(n813) );
  NAND2X2 U1794 ( .A(\sigadd/N22 ), .B(n501), .Y(n814) );
  NAND2X2 U1795 ( .A(\sigadd/N27 ), .B(n501), .Y(n809) );
  NAND2X2 U1796 ( .A(\sigadd/N25 ), .B(n501), .Y(n811) );
  NAND2X2 U1797 ( .A(\sigadd/N26 ), .B(n501), .Y(n810) );
  NAND2X2 U1798 ( .A(\sigadd/N29 ), .B(D[31]), .Y(n807) );
  OAI21X4 U1799 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n602), .B0(n806), .Y(
        add_out[28]) );
  NAND2X2 U1800 ( .A(\sigadd/N30 ), .B(D[31]), .Y(n806) );
  NAND2X2 U1801 ( .A(\sigadd/N32 ), .B(D[31]), .Y(n804) );
  NAND2X2 U1802 ( .A(\sigadd/N28 ), .B(n501), .Y(n808) );
  OAI21X4 U1803 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n611), .B0(n801), .Y(
        add_out[33]) );
  NAND2X2 U1804 ( .A(\sigadd/N35 ), .B(D[31]), .Y(n801) );
  NAND2X2 U1805 ( .A(\sigadd/N33 ), .B(D[31]), .Y(n803) );
  NAND2X2 U1806 ( .A(\sigadd/N34 ), .B(D[31]), .Y(n802) );
  OAI21X4 U1807 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n584), .B0(n800), .Y(
        add_out[34]) );
  NAND2X2 U1808 ( .A(\sigadd/N36 ), .B(D[31]), .Y(n800) );
  OAI21X4 U1809 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n590), .B0(n799), .Y(
        add_out[35]) );
  NAND2X2 U1810 ( .A(\sigadd/N37 ), .B(D[31]), .Y(n799) );
  OAI21X4 U1811 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n583), .B0(n798), .Y(
        \normal/srl_15/A[36] ) );
  NAND2X2 U1812 ( .A(\sigadd/N38 ), .B(D[31]), .Y(n798) );
  NAND2X2 U1813 ( .A(\sigadd/N39 ), .B(D[31]), .Y(n797) );
  OAI21X4 U1814 ( .A0(\sigadd/sub_add_11_b0/B[49] ), .A1(n582), .B0(n796), .Y(
        add_out[38]) );
  NAND2X2 U1815 ( .A(\sigadd/N40 ), .B(D[31]), .Y(n796) );
  NAND2X2 U1816 ( .A(\sigadd/N41 ), .B(D[31]), .Y(n795) );
  NAND2X2 U1817 ( .A(\sigadd/N42 ), .B(D[31]), .Y(n794) );
  INVX2 U1818 ( .A(\sigadd/sig[3] ), .Y(\sigadd/sub_add_11_b0/n96 ) );
  INVX2 U1819 ( .A(\sigadd/sig[4] ), .Y(\sigadd/sub_add_11_b0/n95 ) );
  OR2X2 U1820 ( .A(ali_P[44]), .B(ali_C[44]), .Y(n619) );
  OR2X2 U1821 ( .A(ali_P[42]), .B(ali_C[42]), .Y(n593) );
  OR2X2 U1822 ( .A(ali_P[40]), .B(ali_C[40]), .Y(n594) );
  OR2X2 U1823 ( .A(ali_P[14]), .B(ali_C[14]), .Y(n547) );
  OR2X2 U1824 ( .A(ali_P[12]), .B(ali_C[12]), .Y(n548) );
  OR2X2 U1825 ( .A(ali_P[10]), .B(ali_C[10]), .Y(n549) );
  INVX2 U1826 ( .A(\sigadd/add_9/n217 ), .Y(\sigadd/add_9/n215 ) );
  OR2X2 U1827 ( .A(ali_P[8]), .B(ali_C[8]), .Y(n550) );
  INVX2 U1828 ( .A(\sigadd/add_9/n225 ), .Y(\sigadd/add_9/n223 ) );
  OR2X2 U1829 ( .A(ali_P[6]), .B(ali_C[6]), .Y(n551) );
  INVX2 U1830 ( .A(\sigadd/add_9/n233 ), .Y(\sigadd/add_9/n231 ) );
  OR2X2 U1831 ( .A(ali_P[4]), .B(ali_C[4]), .Y(n552) );
  INVX2 U1832 ( .A(\sigadd/add_9/n241 ), .Y(\sigadd/add_9/n239 ) );
  INVX2 U1833 ( .A(\sigadd/sig[1] ), .Y(\sigadd/sub_add_11_b0/n98 ) );
  INVX2 U1834 ( .A(\sigadd/sig[2] ), .Y(\sigadd/sub_add_11_b0/n97 ) );
  OR2X2 U1835 ( .A(ali_P[2]), .B(ali_C[2]), .Y(n553) );
  INVX2 U1836 ( .A(\mul/mult_6/n125 ), .Y(sig_P[0]) );
  NAND2BX2 U1837 ( .AN(\selc/N209 ), .B(\two_en[1] ), .Y(sel_C[46]) );
  INVX2 U1838 ( .A(sig_C[45]), .Y(\selc/r300/A[45] ) );
  INVX2 U1839 ( .A(sig_C[44]), .Y(\selc/r300/A[44] ) );
  INVX2 U1840 ( .A(sig_C[43]), .Y(\selc/r300/A[43] ) );
  INVX2 U1841 ( .A(sig_C[42]), .Y(\selc/r300/A[42] ) );
  INVX2 U1842 ( .A(sig_C[41]), .Y(\selc/r300/A[41] ) );
  INVX2 U1843 ( .A(sig_C[40]), .Y(\selc/r300/A[40] ) );
  INVX2 U1844 ( .A(sig_C[39]), .Y(\selc/r300/A[39] ) );
  INVX2 U1845 ( .A(sig_C[38]), .Y(\selc/r300/A[38] ) );
  INVX2 U1846 ( .A(sig_C[37]), .Y(\selc/r300/A[37] ) );
  INVX2 U1847 ( .A(sig_C[36]), .Y(\selc/r300/A[36] ) );
  INVX2 U1848 ( .A(sig_C[35]), .Y(\selc/r300/A[35] ) );
  INVX2 U1849 ( .A(sig_C[34]), .Y(\selc/r300/A[34] ) );
  INVX2 U1850 ( .A(sig_C[33]), .Y(\selc/r300/A[33] ) );
  INVX2 U1851 ( .A(sig_C[32]), .Y(\selc/r300/A[32] ) );
  INVX2 U1852 ( .A(sig_C[31]), .Y(\selc/r300/A[31] ) );
  INVX2 U1853 ( .A(sig_C[30]), .Y(\selc/r300/A[30] ) );
  INVX2 U1854 ( .A(sig_C[29]), .Y(\selc/r300/A[29] ) );
  INVX2 U1855 ( .A(sig_C[28]), .Y(\selc/r300/A[28] ) );
  INVX2 U1856 ( .A(sig_C[27]), .Y(\selc/r300/A[27] ) );
  INVX2 U1857 ( .A(sig_C[26]), .Y(\selc/r300/A[26] ) );
  INVX2 U1858 ( .A(sig_C[25]), .Y(\selc/r300/A[25] ) );
  INVX2 U1859 ( .A(sig_C[24]), .Y(\selc/r300/A[24] ) );
  INVX4 U1860 ( .A(\two_en[1] ), .Y(n720) );
  NAND2X2 U1861 ( .A(\selc/N161 ), .B(n502), .Y(n727) );
  NAND2X2 U1862 ( .A(\selc/N160 ), .B(n502), .Y(n728) );
  NAND2X2 U1863 ( .A(\selc/N159 ), .B(n502), .Y(n729) );
  NAND2X2 U1864 ( .A(\selc/N158 ), .B(n502), .Y(n730) );
  NAND2X2 U1865 ( .A(\selc/N157 ), .B(n724), .Y(n731) );
  NAND2X2 U1866 ( .A(\selc/N156 ), .B(n724), .Y(n732) );
  NAND2X2 U1867 ( .A(\selc/N155 ), .B(n724), .Y(n733) );
  NAND2X2 U1868 ( .A(\selc/N154 ), .B(n502), .Y(n734) );
  NAND2X2 U1869 ( .A(\selc/N153 ), .B(n724), .Y(n735) );
  NAND2X2 U1870 ( .A(\selc/N152 ), .B(n724), .Y(n736) );
  NAND2X2 U1871 ( .A(\selc/N151 ), .B(n502), .Y(n737) );
  NAND2X2 U1872 ( .A(\selc/N150 ), .B(n502), .Y(n738) );
  NAND2X2 U1873 ( .A(\selc/N149 ), .B(n502), .Y(n739) );
  NAND2X2 U1874 ( .A(\selc/N148 ), .B(n502), .Y(n740) );
  OR2X2 U1875 ( .A(sub_out[6]), .B(sub_out[7]), .Y(\align/sra_10/n254 ) );
  INVX2 U1876 ( .A(exp_C[0]), .Y(\sub/r301/n17 ) );
  INVX2 U1877 ( .A(exp_C[4]), .Y(\sub/r301/n13 ) );
  INVX2 U1878 ( .A(exp_P[2]), .Y(\sub/sub_17/n15 ) );
  INVX2 U1879 ( .A(exp_P[3]), .Y(\sub/sub_17/n14 ) );
  INVX2 U1880 ( .A(sig_P[40]), .Y(\selc/r299/A[40] ) );
  INVX2 U1881 ( .A(sig_P[39]), .Y(\selc/r299/A[39] ) );
  INVX2 U1882 ( .A(sig_P[38]), .Y(\selc/r299/A[38] ) );
  INVX2 U1883 ( .A(sig_P[37]), .Y(\selc/r299/A[37] ) );
  INVX2 U1884 ( .A(sig_P[36]), .Y(\selc/r299/A[36] ) );
  INVX2 U1885 ( .A(sig_P[35]), .Y(\selc/r299/A[35] ) );
  INVX2 U1886 ( .A(sig_P[34]), .Y(\selc/r299/A[34] ) );
  INVX2 U1887 ( .A(sig_P[33]), .Y(\selc/r299/A[33] ) );
  INVX2 U1888 ( .A(sig_P[32]), .Y(\selc/r299/A[32] ) );
  INVX2 U1889 ( .A(sig_P[31]), .Y(\selc/r299/A[31] ) );
  INVX2 U1890 ( .A(sig_P[30]), .Y(\selc/r299/A[30] ) );
  INVX2 U1891 ( .A(sig_P[29]), .Y(\selc/r299/A[29] ) );
  INVX2 U1892 ( .A(sig_P[28]), .Y(\selc/r299/A[28] ) );
  INVX2 U1893 ( .A(sig_P[27]), .Y(\selc/r299/A[27] ) );
  INVX2 U1894 ( .A(sig_P[26]), .Y(\selc/r299/A[26] ) );
  INVX2 U1895 ( .A(sig_P[25]), .Y(\selc/r299/A[25] ) );
  INVX2 U1896 ( .A(sig_P[24]), .Y(\selc/r299/A[24] ) );
  INVX2 U1897 ( .A(sig_P[23]), .Y(\selc/r299/A[23] ) );
  INVX2 U1898 ( .A(sig_P[22]), .Y(\selc/r299/A[22] ) );
  INVX2 U1899 ( .A(sig_P[21]), .Y(\selc/r299/A[21] ) );
  INVX2 U1900 ( .A(sig_P[20]), .Y(\selc/r299/A[20] ) );
  INVX2 U1901 ( .A(sig_P[19]), .Y(\selc/r299/A[19] ) );
  INVX2 U1902 ( .A(sig_P[18]), .Y(\selc/r299/A[18] ) );
  INVX2 U1903 ( .A(sig_P[17]), .Y(\selc/r299/A[17] ) );
  INVX2 U1904 ( .A(sig_P[16]), .Y(\selc/r299/A[16] ) );
  INVX2 U1905 ( .A(sig_P[15]), .Y(\selc/r299/A[15] ) );
  INVX2 U1906 ( .A(sig_P[14]), .Y(\selc/r299/A[14] ) );
  INVX2 U1907 ( .A(sig_P[13]), .Y(\selc/r299/A[13] ) );
  INVX2 U1908 ( .A(sig_P[12]), .Y(\selc/r299/A[12] ) );
  INVX2 U1909 ( .A(sig_P[11]), .Y(\selc/r299/A[11] ) );
  INVX2 U1910 ( .A(sig_P[10]), .Y(\selc/r299/A[10] ) );
  INVX2 U1911 ( .A(sig_P[9]), .Y(\selc/r299/A[9] ) );
  INVX2 U1912 ( .A(sig_P[8]), .Y(\selc/r299/A[8] ) );
  INVX2 U1913 ( .A(sig_P[7]), .Y(\selc/r299/A[7] ) );
  INVX2 U1914 ( .A(sig_P[6]), .Y(\selc/r299/A[6] ) );
  INVX2 U1915 ( .A(sig_P[5]), .Y(\selc/r299/A[5] ) );
  INVX2 U1916 ( .A(sig_P[4]), .Y(\selc/r299/A[4] ) );
  INVX2 U1917 ( .A(sig_P[3]), .Y(\selc/r299/A[3] ) );
  INVX2 U1918 ( .A(sig_P[2]), .Y(\selc/r299/A[2] ) );
  INVX2 U1919 ( .A(\mul/mult_6/n702 ), .Y(\mul/mult_6/n730 ) );
  INVX2 U1920 ( .A(\mul/mult_6/n675 ), .Y(\mul/mult_6/n725 ) );
  INVX2 U1921 ( .A(\mul/mult_6/n78 ), .Y(n697) );
  INVX2 U1922 ( .A(\mul/mult_6/n587 ), .Y(\mul/mult_6/n585 ) );
  INVX2 U1923 ( .A(sig_P[1]), .Y(\selc/r299/A[1] ) );
  OR2X2 U1924 ( .A(sig_B[0]), .B(sig_B[1]), .Y(n562) );
  NAND2X2 U1925 ( .A(n781), .B(n780), .Y(n783) );
  NAND2X2 U1926 ( .A(n778), .B(n1051), .Y(n779) );
  INVX2 U1927 ( .A(exp_P[1]), .Y(n1045) );
  INVX2 U1928 ( .A(exp_P[5]), .Y(n1047) );
  NOR2X2 U1929 ( .A(n1052), .B(n776), .Y(n777) );
  INVX2 U1930 ( .A(exp_C[1]), .Y(n1028) );
  INVX2 U1931 ( .A(exp_C[2]), .Y(n1061) );
  INVX2 U1932 ( .A(\expadd/add_0_root_sub_0_root_sub_8/n2 ), .Y(exp_P[0]) );
  OR2X2 U1933 ( .A(\expadd/add_0_root_sub_0_root_sub_8/B[0] ), .B(exp_B[0]), 
        .Y(n657) );
  NAND2BX2 U1934 ( .AN(exp_P[4]), .B(exp_C[4]), .Y(n726) );
  INVX2 U1935 ( .A(exp_C[3]), .Y(n1049) );
  INVX2 U1936 ( .A(exp_C[5]), .Y(n1029) );
  INVX2 U1937 ( .A(exp_C[6]), .Y(n1032) );
  INVX2 U1938 ( .A(exp_P[4]), .Y(n1046) );
  INVX2 U1939 ( .A(\expadd/add_0_root_sub_0_root_sub_8/n11 ), .Y(
        \expadd/add_0_root_sub_0_root_sub_8/n9 ) );
  MXI2X1 U1940 ( .A(n1032), .B(n1031), .S0(n516), .Y(
        \ctrl/add_1_root_add_16_2/n13 ) );
  MXI2X1 U1941 ( .A(n1061), .B(\sub/sub_17/n15 ), .S0(n516), .Y(
        \ctrl/add_1_root_add_16_2/A[2] ) );
  OAI21X1 U1942 ( .A0(n1043), .A1(n974), .B0(n973), .Y(n975) );
  AOI21X1 U1943 ( .A0(n972), .A1(add_out[47]), .B0(add_out[49]), .Y(n973) );
  AOI21X1 U1944 ( .A0(n971), .A1(add_out[43]), .B0(add_out[45]), .Y(n974) );
  OAI21X1 U1945 ( .A0(n970), .A1(add_out[28]), .B0(n969), .Y(n976) );
  OAI31X1 U1946 ( .A0(n941), .A1(n927), .A2(n952), .B0(n926), .Y(n928) );
  OAI22X1 U1947 ( .A0(n913), .A1(n912), .B0(n911), .B1(n910), .Y(n914) );
  AOI21X1 U1948 ( .A0(n908), .A1(add_out[39]), .B0(\normal/srl_15/A[41] ), .Y(
        n911) );
  AOI21X1 U1949 ( .A0(n907), .A1(add_out[23]), .B0(\normal/srl_15/A[25] ), .Y(
        n912) );
  OAI22X1 U1950 ( .A0(n890), .A1(n889), .B0(n888), .B1(n897), .Y(n891) );
  NOR3X1 U1951 ( .A(add_out[38]), .B(\normal/srl_15/A[36] ), .C(add_out[34]), 
        .Y(n888) );
  AOI21X1 U1952 ( .A0(n884), .A1(add_out[31]), .B0(add_out[33]), .Y(n886) );
  OAI211XL U1953 ( .A0(n949), .A1(n948), .B0(n947), .C0(n946), .Y(n950) );
  NAND3XL U1954 ( .A(n999), .B(n945), .C(n944), .Y(n946) );
  NOR2XL U1955 ( .A(add_out[48]), .B(add_out[49]), .Y(n947) );
  NOR3BX1 U1956 ( .AN(n943), .B(n942), .C(add_out[33]), .Y(n951) );
  NOR3X1 U1957 ( .A(n940), .B(n939), .C(add_out[17]), .Y(n960) );
  NOR3X1 U1958 ( .A(n968), .B(n938), .C(add_out[13]), .Y(n961) );
  OAI21X1 U1959 ( .A0(\normal/srl_15/A[22] ), .A1(\normal/srl_15/A[25] ), .B0(
        n930), .Y(n876) );
  OAI22X1 U1960 ( .A0(n964), .A1(n862), .B0(n861), .B1(n860), .Y(n863) );
  AOI31X1 U1961 ( .A0(n866), .A1(n851), .A2(\sigadd/sig[0] ), .B0(n850), .Y(
        n857) );
  XNOR2X1 U1962 ( .A(\sigadd/add_9/n229 ), .B(\sigadd/add_9/n45 ), .Y(n656) );
  XOR2X1 U1963 ( .A(\sigadd/add_9/n226 ), .B(\sigadd/add_9/n44 ), .Y(n649) );
  XNOR2X1 U1964 ( .A(\sigadd/add_9/n221 ), .B(\sigadd/add_9/n43 ), .Y(n648) );
  XOR2X1 U1965 ( .A(\sigadd/add_9/n218 ), .B(\sigadd/add_9/n42 ), .Y(n636) );
  XNOR2X1 U1966 ( .A(\sigadd/add_9/n213 ), .B(\sigadd/add_9/n41 ), .Y(n647) );
  XOR2X1 U1967 ( .A(\sigadd/add_9/n210 ), .B(\sigadd/add_9/n40 ), .Y(n635) );
  XNOR2X1 U1968 ( .A(\sigadd/add_9/n205 ), .B(\sigadd/add_9/n39 ), .Y(n646) );
  XOR2X1 U1969 ( .A(\sigadd/add_9/n202 ), .B(\sigadd/add_9/n38 ), .Y(n634) );
  XNOR2X1 U1970 ( .A(\sigadd/add_9/n197 ), .B(\sigadd/add_9/n37 ), .Y(n645) );
  XOR2X1 U1971 ( .A(\sigadd/add_9/n194 ), .B(\sigadd/add_9/n36 ), .Y(n633) );
  XNOR2X1 U1972 ( .A(\sigadd/add_9/n189 ), .B(\sigadd/add_9/n35 ), .Y(n644) );
  XOR2X1 U1973 ( .A(\sigadd/add_9/n186 ), .B(\sigadd/add_9/n34 ), .Y(n623) );
  XNOR2X1 U1974 ( .A(\sigadd/add_9/n181 ), .B(\sigadd/add_9/n33 ), .Y(n632) );
  XOR2X1 U1975 ( .A(\sigadd/add_9/n178 ), .B(\sigadd/add_9/n32 ), .Y(n622) );
  XNOR2X1 U1976 ( .A(\sigadd/add_9/n173 ), .B(\sigadd/add_9/n31 ), .Y(n631) );
  XOR2X1 U1977 ( .A(\sigadd/add_9/n170 ), .B(\sigadd/add_9/n30 ), .Y(n621) );
  XNOR2X1 U1978 ( .A(\sigadd/add_9/n165 ), .B(\sigadd/add_9/n29 ), .Y(n630) );
  XOR2X1 U1979 ( .A(\sigadd/add_9/n162 ), .B(\sigadd/add_9/n28 ), .Y(n620) );
  XNOR2X1 U1980 ( .A(\sigadd/add_9/n157 ), .B(\sigadd/add_9/n27 ), .Y(n616) );
  XOR2X1 U1981 ( .A(\sigadd/add_9/n154 ), .B(\sigadd/add_9/n26 ), .Y(n604) );
  XNOR2X1 U1982 ( .A(\sigadd/add_9/n149 ), .B(\sigadd/add_9/n25 ), .Y(n615) );
  XOR2X1 U1983 ( .A(\sigadd/add_9/n146 ), .B(\sigadd/add_9/n24 ), .Y(n603) );
  XNOR2X1 U1984 ( .A(\sigadd/add_9/n141 ), .B(\sigadd/add_9/n23 ), .Y(n614) );
  XOR2X1 U1985 ( .A(\sigadd/add_9/n138 ), .B(\sigadd/add_9/n22 ), .Y(n602) );
  XNOR2X1 U1986 ( .A(\sigadd/add_9/n133 ), .B(\sigadd/add_9/n21 ), .Y(n613) );
  XOR2X1 U1987 ( .A(\sigadd/add_9/n130 ), .B(\sigadd/add_9/n20 ), .Y(n601) );
  XNOR2X1 U1988 ( .A(\sigadd/add_9/n125 ), .B(\sigadd/add_9/n19 ), .Y(n612) );
  XOR2X1 U1989 ( .A(\sigadd/add_9/n122 ), .B(\sigadd/add_9/n18 ), .Y(n600) );
  XNOR2X1 U1990 ( .A(\sigadd/add_9/n117 ), .B(\sigadd/add_9/n17 ), .Y(n611) );
  XOR2X1 U1991 ( .A(\sigadd/add_9/n114 ), .B(\sigadd/add_9/n16 ), .Y(n584) );
  XNOR2X1 U1992 ( .A(\sigadd/add_9/n77 ), .B(\sigadd/add_9/n7 ), .Y(n567) );
  MX2X1 U1993 ( .A(\align/N100 ), .B(sel_C[46]), .S0(n787), .Y(ali_C[46]) );
  MX2X1 U1994 ( .A(\align/N99 ), .B(sel_C[45]), .S0(n787), .Y(ali_C[45]) );
  MX2X1 U1995 ( .A(\align/N98 ), .B(sel_C[44]), .S0(n787), .Y(ali_C[44]) );
  MX2X1 U1996 ( .A(\align/N97 ), .B(sel_C[43]), .S0(n787), .Y(ali_C[43]) );
  MX2X1 U1997 ( .A(\align/N96 ), .B(sel_C[42]), .S0(n787), .Y(ali_C[42]) );
  MX2X1 U1998 ( .A(\align/N95 ), .B(sel_C[41]), .S0(n787), .Y(ali_C[41]) );
  MX2X1 U1999 ( .A(\align/N94 ), .B(sel_C[40]), .S0(n787), .Y(ali_C[40]) );
  MX2X1 U2000 ( .A(\align/N93 ), .B(sel_C[39]), .S0(n787), .Y(ali_C[39]) );
  MX2X1 U2001 ( .A(\align/N92 ), .B(sel_C[38]), .S0(n787), .Y(ali_C[38]) );
  MX2X1 U2002 ( .A(\align/N91 ), .B(sel_C[37]), .S0(n787), .Y(ali_C[37]) );
  MX2X1 U2003 ( .A(\align/N90 ), .B(sel_C[36]), .S0(n787), .Y(ali_C[36]) );
  MX2X1 U2004 ( .A(\align/N89 ), .B(sel_C[35]), .S0(n787), .Y(ali_C[35]) );
  MX2X1 U2005 ( .A(\align/N88 ), .B(sel_C[34]), .S0(n787), .Y(ali_C[34]) );
  MX2X1 U2006 ( .A(\align/N87 ), .B(sel_C[33]), .S0(n787), .Y(ali_C[33]) );
  MX2X1 U2007 ( .A(\align/N86 ), .B(sel_C[32]), .S0(n787), .Y(ali_C[32]) );
  MX2X1 U2008 ( .A(\align/N85 ), .B(sel_C[31]), .S0(n787), .Y(ali_C[31]) );
  MX2X1 U2009 ( .A(\align/N84 ), .B(sel_C[30]), .S0(n787), .Y(ali_C[30]) );
  MX2X1 U2010 ( .A(\align/N83 ), .B(sel_C[29]), .S0(n787), .Y(ali_C[29]) );
  MX2X1 U2011 ( .A(\align/N82 ), .B(sel_C[28]), .S0(n787), .Y(ali_C[28]) );
  MX2X1 U2012 ( .A(\align/N81 ), .B(sel_C[27]), .S0(n787), .Y(ali_C[27]) );
  MX2X1 U2013 ( .A(\align/N80 ), .B(sel_C[26]), .S0(n787), .Y(ali_C[26]) );
  MX2X1 U2014 ( .A(\align/N79 ), .B(sel_C[25]), .S0(n787), .Y(ali_C[25]) );
  MX2X1 U2015 ( .A(\align/N78 ), .B(sel_C[24]), .S0(n787), .Y(ali_C[24]) );
  MX2X1 U2016 ( .A(\align/N77 ), .B(sel_C[23]), .S0(n787), .Y(ali_C[23]) );
  NOR2BX1 U2017 ( .AN(\align/N76 ), .B(n787), .Y(ali_C[22]) );
  NOR2BX1 U2018 ( .AN(\align/N75 ), .B(n787), .Y(ali_C[21]) );
  NOR2BX1 U2019 ( .AN(\align/N74 ), .B(n787), .Y(ali_C[20]) );
  NOR2BX1 U2020 ( .AN(\align/N73 ), .B(n787), .Y(ali_C[19]) );
  NOR2BX1 U2021 ( .AN(\align/N72 ), .B(n787), .Y(ali_C[18]) );
  NOR2BX1 U2022 ( .AN(\align/N71 ), .B(n787), .Y(ali_C[17]) );
  NOR2BX1 U2023 ( .AN(\align/N70 ), .B(n787), .Y(ali_C[16]) );
  NOR2BX1 U2024 ( .AN(\align/N69 ), .B(n787), .Y(ali_C[15]) );
  NOR2BX1 U2025 ( .AN(\align/N68 ), .B(n787), .Y(ali_C[14]) );
  NOR2BX1 U2026 ( .AN(\align/N67 ), .B(n787), .Y(ali_C[13]) );
  NOR2BX1 U2027 ( .AN(\align/N66 ), .B(n787), .Y(ali_C[12]) );
  NOR2BX1 U2028 ( .AN(\align/N65 ), .B(n787), .Y(ali_C[11]) );
  NOR2BX1 U2029 ( .AN(\align/N64 ), .B(n787), .Y(ali_C[10]) );
  NOR2BX1 U2030 ( .AN(\align/N63 ), .B(n787), .Y(ali_C[9]) );
  NOR2BX1 U2031 ( .AN(\align/N62 ), .B(n787), .Y(ali_C[8]) );
  NOR2BX1 U2032 ( .AN(\align/N61 ), .B(n787), .Y(ali_C[7]) );
  NOR2BX1 U2033 ( .AN(n719), .B(\align/sra_11/n483 ), .Y(\align/sra_11/n480 )
         );
  NOR2BX1 U2034 ( .AN(\align/N60 ), .B(n787), .Y(ali_C[6]) );
  NOR2BX1 U2035 ( .AN(n719), .B(\align/sra_11/n492 ), .Y(\align/sra_11/n489 )
         );
  NOR2BX1 U2036 ( .AN(\align/N59 ), .B(n787), .Y(ali_C[5]) );
  NOR2BX1 U2037 ( .AN(n719), .B(\align/sra_11/n501 ), .Y(\align/sra_11/n498 )
         );
  NOR2BX1 U2038 ( .AN(\align/N58 ), .B(n787), .Y(ali_C[4]) );
  NOR2BX1 U2039 ( .AN(n719), .B(\align/sra_11/n510 ), .Y(\align/sra_11/n507 )
         );
  NOR2BX1 U2040 ( .AN(\align/N57 ), .B(n787), .Y(ali_C[3]) );
  NOR2BX1 U2041 ( .AN(n719), .B(\align/sra_11/n537 ), .Y(\align/sra_11/n534 )
         );
  NOR2BX1 U2042 ( .AN(n511), .B(\align/sra_11/n677 ), .Y(\align/sra_11/n646 )
         );
  NOR2BX1 U2043 ( .AN(\align/N56 ), .B(n787), .Y(ali_C[2]) );
  NOR2BX1 U2044 ( .AN(n719), .B(\align/sra_11/n573 ), .Y(\align/sra_11/n570 )
         );
  NOR2BX1 U2045 ( .AN(n511), .B(\align/sra_11/n689 ), .Y(\align/sra_11/n652 )
         );
  MX2X1 U2046 ( .A(\align/N6 ), .B(sel_P[2]), .S0(n516), .Y(ali_P[2]) );
  NOR2BX1 U2047 ( .AN(n511), .B(\align/sra_11/n723 ), .Y(\align/sra_11/n478 )
         );
  NOR2BX1 U2048 ( .AN(\align/N55 ), .B(n787), .Y(ali_C[1]) );
  MX2X1 U2049 ( .A(sig_C[45]), .B(\selc/N208 ), .S0(\two_en[1] ), .Y(sel_C[45]) );
  MX2X1 U2050 ( .A(sig_C[44]), .B(\selc/N207 ), .S0(\two_en[1] ), .Y(sel_C[44]) );
  MX2X1 U2051 ( .A(sig_C[43]), .B(\selc/N206 ), .S0(\two_en[1] ), .Y(sel_C[43]) );
  MX2X1 U2052 ( .A(sig_C[42]), .B(\selc/N205 ), .S0(\two_en[1] ), .Y(sel_C[42]) );
  MX2X1 U2053 ( .A(sig_C[41]), .B(\selc/N204 ), .S0(\two_en[1] ), .Y(sel_C[41]) );
  MX2X1 U2054 ( .A(sig_C[40]), .B(\selc/N203 ), .S0(\two_en[1] ), .Y(sel_C[40]) );
  MX2X1 U2055 ( .A(sig_C[39]), .B(\selc/N202 ), .S0(\two_en[1] ), .Y(sel_C[39]) );
  MX2X1 U2056 ( .A(sig_C[38]), .B(\selc/N201 ), .S0(\two_en[1] ), .Y(sel_C[38]) );
  MX2X1 U2057 ( .A(sig_C[37]), .B(\selc/N200 ), .S0(\two_en[1] ), .Y(sel_C[37]) );
  MX2X1 U2058 ( .A(sig_C[36]), .B(\selc/N199 ), .S0(\two_en[1] ), .Y(sel_C[36]) );
  MX2X1 U2059 ( .A(sig_C[35]), .B(\selc/N198 ), .S0(\two_en[1] ), .Y(sel_C[35]) );
  MX2X1 U2060 ( .A(sig_C[34]), .B(\selc/N197 ), .S0(\two_en[1] ), .Y(sel_C[34]) );
  MX2X1 U2061 ( .A(sig_C[33]), .B(\selc/N196 ), .S0(\two_en[1] ), .Y(sel_C[33]) );
  NOR2BX1 U2062 ( .AN(n719), .B(\align/sra_11/n636 ), .Y(\align/sra_11/n633 )
         );
  MX2X1 U2063 ( .A(sig_C[32]), .B(\selc/N195 ), .S0(\two_en[1] ), .Y(sel_C[32]) );
  MX2X1 U2064 ( .A(sig_C[31]), .B(\selc/N194 ), .S0(\two_en[1] ), .Y(sel_C[31]) );
  MX2X1 U2065 ( .A(sig_C[30]), .B(\selc/N193 ), .S0(\two_en[1] ), .Y(sel_C[30]) );
  MX2X1 U2066 ( .A(sig_C[29]), .B(\selc/N192 ), .S0(\two_en[1] ), .Y(sel_C[29]) );
  MX2X1 U2067 ( .A(sig_C[28]), .B(\selc/N191 ), .S0(\two_en[1] ), .Y(sel_C[28]) );
  MX2X1 U2068 ( .A(sig_C[27]), .B(\selc/N190 ), .S0(\two_en[1] ), .Y(sel_C[27]) );
  MX2X1 U2069 ( .A(sig_C[26]), .B(\selc/N189 ), .S0(\two_en[1] ), .Y(sel_C[26]) );
  MX2X1 U2070 ( .A(sig_C[25]), .B(\selc/N188 ), .S0(\two_en[1] ), .Y(sel_C[25]) );
  NOR2BX1 U2071 ( .AN(n511), .B(\align/sra_11/n663 ), .Y(\align/sra_11/n471 )
         );
  MX2X1 U2072 ( .A(sig_C[24]), .B(\selc/N187 ), .S0(\two_en[1] ), .Y(sel_C[24]) );
  MX2X1 U2073 ( .A(sig_C[23]), .B(sig_C[23]), .S0(\two_en[1] ), .Y(sel_C[23])
         );
  MX2X1 U2074 ( .A(\align/N5 ), .B(sel_P[1]), .S0(n516), .Y(ali_P[1]) );
  OAI21X1 U2075 ( .A0(n502), .A1(\selc/r299/A[32] ), .B0(n743), .Y(sel_P[32])
         );
  OAI21X1 U2076 ( .A0(n502), .A1(\selc/r299/A[31] ), .B0(n744), .Y(sel_P[31])
         );
  OAI21X1 U2077 ( .A0(n502), .A1(\selc/r299/A[30] ), .B0(n745), .Y(sel_P[30])
         );
  OAI21X1 U2078 ( .A0(n502), .A1(\selc/r299/A[29] ), .B0(n746), .Y(sel_P[29])
         );
  OAI21X1 U2079 ( .A0(n502), .A1(\selc/r299/A[28] ), .B0(n747), .Y(sel_P[28])
         );
  OAI21X1 U2080 ( .A0(n502), .A1(\selc/r299/A[27] ), .B0(n748), .Y(sel_P[27])
         );
  OAI21X1 U2081 ( .A0(n502), .A1(\selc/r299/A[26] ), .B0(n749), .Y(sel_P[26])
         );
  OAI21X1 U2082 ( .A0(n502), .A1(\selc/r299/A[25] ), .B0(n750), .Y(sel_P[25])
         );
  OAI21X1 U2083 ( .A0(n502), .A1(\selc/r299/A[24] ), .B0(n751), .Y(sel_P[24])
         );
  OAI21X1 U2084 ( .A0(n502), .A1(\selc/r299/A[23] ), .B0(n752), .Y(sel_P[23])
         );
  OAI21X1 U2085 ( .A0(n502), .A1(\selc/r299/A[22] ), .B0(n753), .Y(sel_P[22])
         );
  OAI21X1 U2086 ( .A0(n502), .A1(\selc/r299/A[21] ), .B0(n754), .Y(sel_P[21])
         );
  OAI21X1 U2087 ( .A0(n502), .A1(\selc/r299/A[20] ), .B0(n755), .Y(sel_P[20])
         );
  OAI21X1 U2088 ( .A0(n502), .A1(\selc/r299/A[19] ), .B0(n756), .Y(sel_P[19])
         );
  OAI21X1 U2089 ( .A0(n502), .A1(\selc/r299/A[18] ), .B0(n757), .Y(sel_P[18])
         );
  OAI21X1 U2090 ( .A0(n502), .A1(\selc/r299/A[17] ), .B0(n758), .Y(sel_P[17])
         );
  OAI21X1 U2091 ( .A0(n502), .A1(\selc/r299/A[34] ), .B0(n741), .Y(sel_P[34])
         );
  OAI21X1 U2092 ( .A0(n502), .A1(\selc/r299/A[33] ), .B0(n742), .Y(sel_P[33])
         );
  OAI21X1 U2093 ( .A0(n502), .A1(\selc/r299/A[16] ), .B0(n759), .Y(sel_P[16])
         );
  OAI21X1 U2094 ( .A0(n502), .A1(\selc/r299/A[15] ), .B0(n760), .Y(sel_P[15])
         );
  OAI21X1 U2095 ( .A0(n502), .A1(\selc/r299/A[14] ), .B0(n761), .Y(sel_P[14])
         );
  OAI21X1 U2096 ( .A0(n502), .A1(\selc/r299/A[13] ), .B0(n762), .Y(sel_P[13])
         );
  OAI21X1 U2097 ( .A0(n502), .A1(\selc/r299/A[12] ), .B0(n763), .Y(sel_P[12])
         );
  OAI21X1 U2098 ( .A0(n502), .A1(\selc/r299/A[11] ), .B0(n764), .Y(sel_P[11])
         );
  OAI21X1 U2099 ( .A0(n502), .A1(\selc/r299/A[10] ), .B0(n765), .Y(sel_P[10])
         );
  OAI21X1 U2100 ( .A0(n502), .A1(\selc/r299/A[9] ), .B0(n766), .Y(sel_P[9]) );
  OAI21X1 U2101 ( .A0(n502), .A1(\selc/r299/A[8] ), .B0(n767), .Y(sel_P[8]) );
  OAI21X1 U2102 ( .A0(n502), .A1(\selc/r299/A[7] ), .B0(n768), .Y(sel_P[7]) );
  OAI21X1 U2103 ( .A0(n502), .A1(\selc/r299/A[6] ), .B0(n769), .Y(sel_P[6]) );
  OAI21X1 U2104 ( .A0(n502), .A1(\selc/r299/A[5] ), .B0(n770), .Y(sel_P[5]) );
  MX2X1 U2105 ( .A(\sub/N15 ), .B(\sub/N6 ), .S0(n516), .Y(sub_out[1]) );
  OAI21X1 U2106 ( .A0(n502), .A1(\selc/r299/A[4] ), .B0(n771), .Y(sel_P[4]) );
  OAI21X1 U2107 ( .A0(n502), .A1(\selc/r299/A[3] ), .B0(n772), .Y(sel_P[3]) );
  OAI21X1 U2108 ( .A0(n502), .A1(\selc/r299/A[2] ), .B0(n773), .Y(sel_P[2]) );
  MX2X1 U2109 ( .A(\sub/N21 ), .B(\sub/N12 ), .S0(n516), .Y(sub_out[7]) );
  MX2X1 U2110 ( .A(\sub/N20 ), .B(\sub/N11 ), .S0(n516), .Y(sub_out[6]) );
  OAI21X1 U2111 ( .A0(n502), .A1(\selc/r299/A[1] ), .B0(n774), .Y(sel_P[1]) );
  MXI2X1 U2112 ( .A(\sub/r301/n13 ), .B(n1046), .S0(n516), .Y(
        \ctrl/add_1_root_add_16_2/A[4] ) );
  OA22X2 U2113 ( .A0(exp_P[2]), .A1(n1061), .B0(exp_P[1]), .B1(n1028), .Y(
        n1044) );
  AOI2BB1X2 U2114 ( .A0N(exp_A[0]), .A1N(exp_A[1]), .B0(n1053), .Y(\expadd/N1 ) );
  CMPR42X1 U2115 ( .A(\mul/mult_6/n472 ), .B(\mul/mult_6/n888 ), .C(
        \mul/mult_6/n473 ), .D(\mul/mult_6/n936 ), .ICI(\mul/mult_6/n912 ), 
        .S(\mul/mult_6/n470 ), .ICO(\mul/mult_6/n468 ), .CO(\mul/mult_6/n469 )
         );
  CMPR42X1 U2116 ( .A(\mul/mult_6/n477 ), .B(\mul/mult_6/n889 ), .C(
        \mul/mult_6/n480 ), .D(\mul/mult_6/n913 ), .ICI(\mul/mult_6/n937 ), 
        .S(\mul/mult_6/n475 ), .ICO(\mul/mult_6/n473 ), .CO(\mul/mult_6/n474 )
         );
  CMPR42X1 U2117 ( .A(\mul/mult_6/n467 ), .B(\mul/mult_6/n911 ), .C(
        \mul/mult_6/n887 ), .D(\mul/mult_6/n468 ), .ICI(\mul/mult_6/n935 ), 
        .S(\mul/mult_6/n465 ), .ICO(\mul/mult_6/n463 ), .CO(\mul/mult_6/n464 )
         );
  CMPR42X1 U2118 ( .A(\mul/mult_6/n425 ), .B(\mul/mult_6/n857 ), .C(
        \mul/mult_6/n833 ), .D(\mul/mult_6/n429 ), .ICI(\mul/mult_6/n905 ), 
        .S(\mul/mult_6/n423 ), .ICO(\mul/mult_6/n421 ), .CO(\mul/mult_6/n422 )
         );
  CMPR42X1 U2119 ( .A(\mul/mult_6/n404 ), .B(\mul/mult_6/n878 ), .C(
        \mul/mult_6/n395 ), .D(\mul/mult_6/n926 ), .ICI(\mul/mult_6/n401 ), 
        .S(\mul/mult_6/n393 ), .ICO(\mul/mult_6/n391 ), .CO(\mul/mult_6/n392 )
         );
  CMPR42X1 U2120 ( .A(\mul/mult_6/n415 ), .B(\mul/mult_6/n832 ), .C(
        \mul/mult_6/n856 ), .D(\mul/mult_6/n880 ), .ICI(\mul/mult_6/n421 ), 
        .S(\mul/mult_6/n413 ), .ICO(\mul/mult_6/n411 ), .CO(\mul/mult_6/n412 )
         );
  CMPR42X1 U2121 ( .A(\mul/mult_6/n441 ), .B(\mul/mult_6/n835 ), .C(
        \mul/mult_6/n447 ), .D(\mul/mult_6/n859 ), .ICI(\mul/mult_6/n907 ), 
        .S(\mul/mult_6/n439 ), .ICO(\mul/mult_6/n437 ), .CO(\mul/mult_6/n438 )
         );
  CMPR42X1 U2122 ( .A(\mul/mult_6/n854 ), .B(\mul/mult_6/n902 ), .C(
        \mul/mult_6/n402 ), .D(\mul/mult_6/n393 ), .ICI(\mul/mult_6/n398 ), 
        .S(\mul/mult_6/n390 ), .ICO(\mul/mult_6/n388 ), .CO(\mul/mult_6/n389 )
         );
  CMPR42X1 U2123 ( .A(\mul/mult_6/n879 ), .B(\mul/mult_6/n927 ), .C(
        \mul/mult_6/n412 ), .D(\mul/mult_6/n403 ), .ICI(\mul/mult_6/n408 ), 
        .S(\mul/mult_6/n400 ), .ICO(\mul/mult_6/n398 ), .CO(\mul/mult_6/n399 )
         );
  CMPR42X1 U2124 ( .A(\mul/mult_6/n881 ), .B(\mul/mult_6/n929 ), .C(
        \mul/mult_6/n430 ), .D(\mul/mult_6/n423 ), .ICI(\mul/mult_6/n426 ), 
        .S(\mul/mult_6/n420 ), .ICO(\mul/mult_6/n418 ), .CO(\mul/mult_6/n419 )
         );
  CMPR42X1 U2125 ( .A(\mul/mult_6/n930 ), .B(\mul/mult_6/n906 ), .C(
        \mul/mult_6/n438 ), .D(\mul/mult_6/n434 ), .ICI(\mul/mult_6/n431 ), 
        .S(\mul/mult_6/n428 ), .ICO(\mul/mult_6/n426 ), .CO(\mul/mult_6/n427 )
         );
  CMPR42X1 U2126 ( .A(\mul/mult_6/n452 ), .B(\mul/mult_6/n932 ), .C(
        \mul/mult_6/n446 ), .D(\mul/mult_6/n908 ), .ICI(\mul/mult_6/n449 ), 
        .S(\mul/mult_6/n444 ), .ICO(\mul/mult_6/n442 ), .CO(\mul/mult_6/n443 )
         );
  CMPR42X1 U2127 ( .A(\mul/mult_6/n883 ), .B(\mul/mult_6/n445 ), .C(
        \mul/mult_6/n931 ), .D(\mul/mult_6/n439 ), .ICI(\mul/mult_6/n442 ), 
        .S(\mul/mult_6/n436 ), .ICO(\mul/mult_6/n434 ), .CO(\mul/mult_6/n435 )
         );
  CMPR42X1 U2128 ( .A(\mul/mult_6/n460 ), .B(\mul/mult_6/n886 ), .C(
        \mul/mult_6/n934 ), .D(\mul/mult_6/n910 ), .ICI(\mul/mult_6/n463 ), 
        .S(\mul/mult_6/n458 ), .ICO(\mul/mult_6/n456 ), .CO(\mul/mult_6/n457 )
         );
  CMPR42X1 U2129 ( .A(\mul/mult_6/n453 ), .B(\mul/mult_6/n909 ), .C(
        \mul/mult_6/n885 ), .D(\mul/mult_6/n933 ), .ICI(\mul/mult_6/n456 ), 
        .S(\mul/mult_6/n451 ), .ICO(\mul/mult_6/n449 ), .CO(\mul/mult_6/n450 )
         );
  CMPR42X1 U2130 ( .A(\mul/mult_6/n433 ), .B(\mul/mult_6/n834 ), .C(
        \mul/mult_6/n437 ), .D(\mul/mult_6/n882 ), .ICI(\mul/mult_6/n858 ), 
        .S(\mul/mult_6/n431 ), .ICO(\mul/mult_6/n429 ), .CO(\mul/mult_6/n430 )
         );
  CMPR42X1 U2131 ( .A(\mul/mult_6/n354 ), .B(\mul/mult_6/n778 ), .C(
        \mul/mult_6/n802 ), .D(\mul/mult_6/n826 ), .ICI(\mul/mult_6/n361 ), 
        .S(\mul/mult_6/n352 ), .ICO(\mul/mult_6/n350 ), .CO(\mul/mult_6/n351 )
         );
  CMPR42X1 U2132 ( .A(\mul/mult_6/n365 ), .B(\mul/mult_6/n803 ), .C(
        \mul/mult_6/n779 ), .D(\mul/mult_6/n372 ), .ICI(\mul/mult_6/n851 ), 
        .S(\mul/mult_6/n363 ), .ICO(\mul/mult_6/n361 ), .CO(\mul/mult_6/n362 )
         );
  CMPR42X1 U2133 ( .A(\mul/mult_6/n800 ), .B(\mul/mult_6/n896 ), .C(
        \mul/mult_6/n848 ), .D(\mul/mult_6/n339 ), .ICI(\mul/mult_6/n336 ), 
        .S(\mul/mult_6/n327 ), .ICO(\mul/mult_6/n325 ), .CO(\mul/mult_6/n326 )
         );
  CMPR42X1 U2134 ( .A(\mul/mult_6/n899 ), .B(\mul/mult_6/n923 ), .C(
        \mul/mult_6/n875 ), .D(\mul/mult_6/n373 ), .ICI(\mul/mult_6/n369 ), 
        .S(\mul/mult_6/n360 ), .ICO(\mul/mult_6/n358 ), .CO(\mul/mult_6/n359 )
         );
  CMPR42X1 U2135 ( .A(\mul/mult_6/n853 ), .B(\mul/mult_6/n394 ), .C(
        \mul/mult_6/n901 ), .D(\mul/mult_6/n877 ), .ICI(\mul/mult_6/n925 ), 
        .S(\mul/mult_6/n382 ), .ICO(\mul/mult_6/n380 ), .CO(\mul/mult_6/n381 )
         );
  CMPR42X1 U2136 ( .A(\mul/mult_6/n825 ), .B(\mul/mult_6/n350 ), .C(
        \mul/mult_6/n873 ), .D(\mul/mult_6/n897 ), .ICI(\mul/mult_6/n341 ), 
        .S(\mul/mult_6/n338 ), .ICO(\mul/mult_6/n336 ), .CO(\mul/mult_6/n337 )
         );
  CMPR42X1 U2137 ( .A(\mul/mult_6/n330 ), .B(\mul/mult_6/n340 ), .C(
        \mul/mult_6/n327 ), .D(\mul/mult_6/n337 ), .ICI(\mul/mult_6/n333 ), 
        .S(\mul/mult_6/n324 ), .ICO(\mul/mult_6/n322 ), .CO(\mul/mult_6/n323 )
         );
  CMPR42X1 U2138 ( .A(\mul/mult_6/n347 ), .B(\mul/mult_6/n351 ), .C(
        \mul/mult_6/n348 ), .D(\mul/mult_6/n338 ), .ICI(\mul/mult_6/n344 ), 
        .S(\mul/mult_6/n335 ), .ICO(\mul/mult_6/n333 ), .CO(\mul/mult_6/n334 )
         );
  CMPR42X1 U2139 ( .A(\mul/mult_6/n827 ), .B(\mul/mult_6/n363 ), .C(
        \mul/mult_6/n370 ), .D(\mul/mult_6/n360 ), .ICI(\mul/mult_6/n366 ), 
        .S(\mul/mult_6/n357 ), .ICO(\mul/mult_6/n355 ), .CO(\mul/mult_6/n356 )
         );
  CMPR42X1 U2140 ( .A(\mul/mult_6/n900 ), .B(\mul/mult_6/n374 ), .C(
        \mul/mult_6/n381 ), .D(\mul/mult_6/n377 ), .ICI(\mul/mult_6/n371 ), 
        .S(\mul/mult_6/n368 ), .ICO(\mul/mult_6/n366 ), .CO(\mul/mult_6/n367 )
         );
  CMPR42X1 U2141 ( .A(\mul/mult_6/n343 ), .B(\mul/mult_6/n801 ), .C(
        \mul/mult_6/n777 ), .D(\mul/mult_6/n849 ), .ICI(\mul/mult_6/n921 ), 
        .S(\mul/mult_6/n341 ), .ICO(\mul/mult_6/n339 ), .CO(\mul/mult_6/n340 )
         );
  CMPR42X1 U2142 ( .A(\mul/mult_6/n331 ), .B(\mul/mult_6/n321 ), .C(
        \mul/mult_6/n775 ), .D(\mul/mult_6/n895 ), .ICI(\mul/mult_6/n823 ), 
        .S(\mul/mult_6/n319 ), .ICO(\mul/mult_6/n317 ), .CO(\mul/mult_6/n318 )
         );
  CMPR42X1 U2143 ( .A(n677), .B(\mul/mult_6/n298 ), .C(n627), .D(
        \mul/mult_6/n772 ), .ICI(\mul/mult_6/n868 ), .S(\mul/mult_6/n287 ), 
        .ICO(\mul/mult_6/n285 ), .CO(\mul/mult_6/n286 ) );
  CMPR42X1 U2144 ( .A(n625), .B(\mul/mult_6/n774 ), .C(\mul/mult_6/n822 ), .D(
        \mul/mult_6/n310 ), .ICI(\mul/mult_6/n317 ), .S(\mul/mult_6/n308 ), 
        .ICO(\mul/mult_6/n306 ), .CO(\mul/mult_6/n307 ) );
  CMPR42X1 U2145 ( .A(\mul/mult_6/n299 ), .B(n624), .C(\mul/mult_6/n797 ), .D(
        \mul/mult_6/n309 ), .ICI(\mul/mult_6/n845 ), .S(\mul/mult_6/n297 ), 
        .ICO(\mul/mult_6/n295 ), .CO(\mul/mult_6/n296 ) );
  CMPR42X1 U2146 ( .A(\mul/mult_6/n773 ), .B(\mul/mult_6/n869 ), .C(
        \mul/mult_6/n821 ), .D(\mul/mult_6/n306 ), .ICI(\mul/mult_6/n303 ), 
        .S(\mul/mult_6/n294 ), .ICO(\mul/mult_6/n292 ), .CO(\mul/mult_6/n293 )
         );
  CMPR42X1 U2147 ( .A(\mul/mult_6/n894 ), .B(\mul/mult_6/n798 ), .C(
        \mul/mult_6/n846 ), .D(\mul/mult_6/n870 ), .ICI(\mul/mult_6/n318 ), 
        .S(\mul/mult_6/n305 ), .ICO(\mul/mult_6/n303 ), .CO(\mul/mult_6/n304 )
         );
  CMPR42X1 U2148 ( .A(\mul/mult_6/n922 ), .B(\mul/mult_6/n874 ), .C(
        \mul/mult_6/n850 ), .D(\mul/mult_6/n898 ), .ICI(\mul/mult_6/n358 ), 
        .S(\mul/mult_6/n349 ), .ICO(\mul/mult_6/n347 ), .CO(\mul/mult_6/n348 )
         );
  CMPR42X1 U2149 ( .A(\mul/mult_6/n286 ), .B(\mul/mult_6/n282 ), .C(
        \mul/mult_6/n283 ), .D(\mul/mult_6/n274 ), .ICI(\mul/mult_6/n279 ), 
        .S(\mul/mult_6/n271 ), .ICO(\mul/mult_6/n269 ), .CO(\mul/mult_6/n270 )
         );
  CMPR42X1 U2150 ( .A(\mul/mult_6/n292 ), .B(\mul/mult_6/n287 ), .C(
        \mul/mult_6/n293 ), .D(\mul/mult_6/n284 ), .ICI(\mul/mult_6/n289 ), 
        .S(\mul/mult_6/n281 ), .ICO(\mul/mult_6/n279 ), .CO(\mul/mult_6/n280 )
         );
  CMPR42X1 U2151 ( .A(\mul/mult_6/n314 ), .B(\mul/mult_6/n308 ), .C(
        \mul/mult_6/n315 ), .D(\mul/mult_6/n305 ), .ICI(\mul/mult_6/n311 ), 
        .S(\mul/mult_6/n302 ), .ICO(\mul/mult_6/n300 ), .CO(\mul/mult_6/n301 )
         );
  CMPR42X1 U2152 ( .A(\mul/mult_6/n325 ), .B(\mul/mult_6/n319 ), .C(
        \mul/mult_6/n326 ), .D(\mul/mult_6/n316 ), .ICI(\mul/mult_6/n322 ), 
        .S(\mul/mult_6/n313 ), .ICO(\mul/mult_6/n311 ), .CO(\mul/mult_6/n312 )
         );
  CMPR42X1 U2153 ( .A(\mul/mult_6/n841 ), .B(\mul/mult_6/n258 ), .C(
        \mul/mult_6/n793 ), .D(\mul/mult_6/n769 ), .ICI(\mul/mult_6/n263 ), 
        .S(\mul/mult_6/n256 ), .ICO(\mul/mult_6/n254 ), .CO(\mul/mult_6/n255 )
         );
  CMPR42X1 U2154 ( .A(\mul/mult_6/n241 ), .B(n637), .C(\mul/mult_6/n248 ), .D(
        \mul/mult_6/n791 ), .ICI(\mul/mult_6/n815 ), .S(\mul/mult_6/n239 ), 
        .ICO(\mul/mult_6/n237 ), .CO(\mul/mult_6/n238 ) );
  CMPR42X1 U2155 ( .A(\mul/mult_6/n237 ), .B(\mul/mult_6/n790 ), .C(
        \mul/mult_6/n232 ), .D(\mul/mult_6/n238 ), .ICI(\mul/mult_6/n234 ), 
        .S(\mul/mult_6/n229 ), .ICO(\mul/mult_6/n227 ), .CO(\mul/mult_6/n228 )
         );
  CMPR42X1 U2156 ( .A(\mul/mult_6/n767 ), .B(\mul/mult_6/n245 ), .C(
        \mul/mult_6/n246 ), .D(\mul/mult_6/n239 ), .ICI(\mul/mult_6/n242 ), 
        .S(\mul/mult_6/n236 ), .ICO(\mul/mult_6/n234 ), .CO(\mul/mult_6/n235 )
         );
  CMPR42X1 U2157 ( .A(\mul/mult_6/n816 ), .B(\mul/mult_6/n792 ), .C(
        \mul/mult_6/n255 ), .D(\mul/mult_6/n247 ), .ICI(\mul/mult_6/n251 ), 
        .S(\mul/mult_6/n244 ), .ICO(\mul/mult_6/n242 ), .CO(\mul/mult_6/n243 )
         );
  CMPR42X1 U2158 ( .A(\mul/mult_6/n276 ), .B(\mul/mult_6/n272 ), .C(
        \mul/mult_6/n265 ), .D(\mul/mult_6/n273 ), .ICI(\mul/mult_6/n269 ), 
        .S(\mul/mult_6/n262 ), .ICO(\mul/mult_6/n260 ), .CO(\mul/mult_6/n261 )
         );
  CMPR42X1 U2159 ( .A(n667), .B(sig_B[7]), .C(sig_B[8]), .D(\mul/mult_6/n770 ), 
        .ICI(n629), .S(\mul/mult_6/n268 ), .ICO(\mul/mult_6/n266 ), .CO(
        \mul/mult_6/n267 ) );
  CMPR42X1 U2160 ( .A(sig_B[6]), .B(n676), .C(n626), .D(\mul/mult_6/n795 ), 
        .ICI(\mul/mult_6/n285 ), .S(\mul/mult_6/n277 ), .ICO(\mul/mult_6/n275 ), .CO(\mul/mult_6/n276 ) );
  CMPR42X1 U2161 ( .A(n665), .B(sig_B[13]), .C(sig_B[14]), .D(n643), .ICI(
        \mul/mult_6/n223 ), .S(\mul/mult_6/n219 ), .ICO(\mul/mult_6/n217 ), 
        .CO(\mul/mult_6/n218 ) );
  CMPR42X1 U2162 ( .A(sig_B[12]), .B(n673), .C(n639), .D(\mul/mult_6/n813 ), 
        .ICI(\mul/mult_6/n230 ), .S(\mul/mult_6/n225 ), .ICO(\mul/mult_6/n223 ), .CO(\mul/mult_6/n224 ) );
  CMPR42X1 U2163 ( .A(\mul/mult_6/n211 ), .B(n651), .C(\mul/mult_6/n206 ), .D(
        \mul/mult_6/n762 ), .ICI(\mul/mult_6/n208 ), .S(\mul/mult_6/n204 ), 
        .ICO(\mul/mult_6/n202 ), .CO(\mul/mult_6/n203 ) );
  CMPR42X1 U2164 ( .A(\mul/mult_6/n787 ), .B(\mul/mult_6/n212 ), .C(
        \mul/mult_6/n763 ), .D(\mul/mult_6/n218 ), .ICI(\mul/mult_6/n214 ), 
        .S(\mul/mult_6/n210 ), .ICO(\mul/mult_6/n208 ), .CO(\mul/mult_6/n209 )
         );
  CMPR42X1 U2165 ( .A(\mul/mult_6/n789 ), .B(\mul/mult_6/n765 ), .C(
        \mul/mult_6/n231 ), .D(\mul/mult_6/n225 ), .ICI(\mul/mult_6/n227 ), 
        .S(\mul/mult_6/n222 ), .ICO(\mul/mult_6/n220 ), .CO(\mul/mult_6/n221 )
         );
  CMPR42X1 U2166 ( .A(n663), .B(sig_B[18]), .C(sig_B[20]), .D(n658), .ICI(
        \mul/mult_6/n189 ), .S(\mul/mult_6/n188 ), .ICO(\mul/mult_6/n186 ), 
        .CO(\mul/mult_6/n187 ) );
  CMPR42X1 U2167 ( .A(n671), .B(\mul/mult_6/n200 ), .C(\mul/mult_6/n760 ), .D(
        n655), .ICI(\mul/mult_6/n197 ), .S(\mul/mult_6/n195 ), .ICO(
        \mul/mult_6/n193 ), .CO(\mul/mult_6/n194 ) );
  CMPR42X1 U2168 ( .A(sig_B[19]), .B(n671), .C(\mul/mult_6/n759 ), .D(n654), 
        .ICI(\mul/mult_6/n193 ), .S(\mul/mult_6/n191 ), .ICO(\mul/mult_6/n189 ), .CO(\mul/mult_6/n190 ) );
  MX2X1 U2169 ( .A(\sub/N14 ), .B(\sub/N5 ), .S0(n516), .Y(sub_out[0]) );
  OAI22X1 U2170 ( .A0(exp_C[1]), .A1(n1045), .B0(exp_C[0]), .B1(
        \expadd/add_0_root_sub_0_root_sub_8/n2 ), .Y(n1048) );
  AOI222XL U2171 ( .A0(n1061), .A1(exp_P[2]), .B0(n1049), .B1(exp_P[3]), .C0(
        n1048), .C1(n1044), .Y(n1050) );
  OAI222X1 U2172 ( .A0(n1047), .A1(exp_C[5]), .B0(n1052), .B1(n1050), .C0(
        n1046), .C1(exp_C[4]), .Y(n1051) );
  AOI21X1 U2173 ( .A0(n1055), .A1(n1054), .B0(n1056), .Y(\expadd/N3 ) );
endmodule

